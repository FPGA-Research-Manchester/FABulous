wire Tile_X9Y1_RES2_I0, Tile_X9Y1_RES2_I1, Tile_X9Y1_RES2_I2, Tile_X9Y1_RES2_I3;
(* keep *) OutPass4_frame_config Tile_X9Y1_E (.I0(Tile_X9Y1_RES2_I0), .I1(Tile_X9Y1_RES2_I1), .I2(Tile_X9Y1_RES2_I2), .I3(Tile_X9Y1_RES2_I3));
endmodule