
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_CLB is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_CLB;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_CLB.all;

entity CLB is

   port( N1BEG : out std_logic_vector (2 downto 0);  N2BEG : out 
         std_logic_vector (5 downto 0);  N4BEG : out std_logic_vector (7 downto
         0);  N1END : in std_logic_vector (2 downto 0);  N2END : in 
         std_logic_vector (5 downto 0);  N4END : in std_logic_vector (7 downto 
         0);  E1BEG : out std_logic_vector (3 downto 0);  E2BEG : out 
         std_logic_vector (7 downto 0);  E1END : in std_logic_vector (3 downto 
         0);  E2END : in std_logic_vector (7 downto 0);  S1BEG : out 
         std_logic_vector (4 downto 0);  S2BEG : out std_logic_vector (9 downto
         0);  S1END : in std_logic_vector (4 downto 0);  S2END : in 
         std_logic_vector (9 downto 0);  W1BEG : out std_logic_vector (5 downto
         0);  W2BEG : out std_logic_vector (11 downto 0);  W1END : in 
         std_logic_vector (5 downto 0);  W2END : in std_logic_vector (11 downto
         0);  MODE, CONFin : in std_logic;  CONFout : out std_logic;  CLK : in 
         std_logic);

end CLB;

architecture SYN_Behavioral of CLB is

   component MUX4D1
      port( I0, I1, I2, I3, S0, S1 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22D1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INVD0
      port( I : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX4ND0
      port( I0, I1, I2, I3, S0, S1 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MAOI22D0
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI221D1
      port( A1, A2, B1, B2, C : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2ND0
      port( I0, I1, S : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI32D1
      port( A1, A2, A3, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211D1
      port( A1, A2, B, C : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21D1
      port( A1, A2, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NR2D0
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CKND2D0
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUFFD16
      port( I : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD16
      port( I : in std_logic;  ZN : out std_logic);
   end component;
   
   component NR2D1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AO22D1
      port( A1, A2, B1, B2 : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2D0
      port( I0, I1, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2D0
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   component INVD1
      port( I : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX4D4
      port( I0, I1, I2, I3, S0, S1 : in std_logic;  Z : out std_logic);
   end component;
   
   component DFQD1
      port( D, CP : in std_logic;  Q : out std_logic);
   end component;
   
   component XOR2D1
      port( A1, A2 : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1282, n1283, n1284, n1285, n1286, n1287, n1291, n1292, n1299, n1300,
      n1301, n1302, n1303, n1304, n1305, n1310, n1311, n1312, n1313, n1314, 
      n1315, n1316, n1317, n1318, n1319, n1325, n1326, n1327, n1328, n1329, 
      n1330, n1331, n1332, n1333, n1334, n1335, n1342, conf_data_2_port, 
      conf_data_1_port, A0, A, AQ, B, BQ, C, CQ, D0, D1, D2, D3, D, DQ, TestIn,
      TestOut, IJ_BEG_12_port, IJ_BEG_11_port, IJ_BEG_10_port, IJ_BEG_9_port, 
      IJ_BEG_8_port, IJ_BEG_7_port, IJ_BEG_6_port, IJ_BEG_5_port, IJ_BEG_4_port
      , IJ_BEG_3_port, IJ_BEG_0_port, OJ_BEG_2_port, OJ_BEG_1_port, 
      OJ_BEG_0_port, Inst_clb_slice_4xLUT4_LUT_D_values_0_port, 
      Inst_clb_slice_4xLUT4_LUT_D_values_1_port, 
      Inst_clb_slice_4xLUT4_LUT_D_values_2_port, 
      Inst_clb_slice_4xLUT4_LUT_D_values_3_port, 
      Inst_clb_slice_4xLUT4_LUT_D_values_4_port, 
      Inst_clb_slice_4xLUT4_LUT_D_values_5_port, 
      Inst_clb_slice_4xLUT4_LUT_D_values_6_port, 
      Inst_clb_slice_4xLUT4_LUT_D_values_7_port, 
      Inst_clb_slice_4xLUT4_LUT_D_values_8_port, 
      Inst_clb_slice_4xLUT4_LUT_D_values_9_port, 
      Inst_clb_slice_4xLUT4_LUT_D_values_10_port, 
      Inst_clb_slice_4xLUT4_LUT_D_values_11_port, 
      Inst_clb_slice_4xLUT4_LUT_D_values_12_port, 
      Inst_clb_slice_4xLUT4_LUT_D_values_13_port, 
      Inst_clb_slice_4xLUT4_LUT_D_values_14_port, 
      Inst_clb_slice_4xLUT4_LUT_C_values_0_port, 
      Inst_clb_slice_4xLUT4_LUT_C_values_1_port, 
      Inst_clb_slice_4xLUT4_LUT_C_values_2_port, 
      Inst_clb_slice_4xLUT4_LUT_C_values_3_port, 
      Inst_clb_slice_4xLUT4_LUT_C_values_4_port, 
      Inst_clb_slice_4xLUT4_LUT_C_values_5_port, 
      Inst_clb_slice_4xLUT4_LUT_C_values_6_port, 
      Inst_clb_slice_4xLUT4_LUT_C_values_7_port, 
      Inst_clb_slice_4xLUT4_LUT_C_values_8_port, 
      Inst_clb_slice_4xLUT4_LUT_C_values_9_port, 
      Inst_clb_slice_4xLUT4_LUT_C_values_10_port, 
      Inst_clb_slice_4xLUT4_LUT_C_values_11_port, 
      Inst_clb_slice_4xLUT4_LUT_C_values_12_port, 
      Inst_clb_slice_4xLUT4_LUT_C_values_13_port, 
      Inst_clb_slice_4xLUT4_LUT_C_values_14_port, 
      Inst_clb_slice_4xLUT4_LUT_C_values_15_port, 
      Inst_clb_slice_4xLUT4_LUT_B_values_0_port, 
      Inst_clb_slice_4xLUT4_LUT_B_values_1_port, 
      Inst_clb_slice_4xLUT4_LUT_B_values_2_port, 
      Inst_clb_slice_4xLUT4_LUT_B_values_3_port, 
      Inst_clb_slice_4xLUT4_LUT_B_values_4_port, 
      Inst_clb_slice_4xLUT4_LUT_B_values_5_port, 
      Inst_clb_slice_4xLUT4_LUT_B_values_6_port, 
      Inst_clb_slice_4xLUT4_LUT_B_values_7_port, 
      Inst_clb_slice_4xLUT4_LUT_B_values_8_port, 
      Inst_clb_slice_4xLUT4_LUT_B_values_9_port, 
      Inst_clb_slice_4xLUT4_LUT_B_values_10_port, 
      Inst_clb_slice_4xLUT4_LUT_B_values_11_port, 
      Inst_clb_slice_4xLUT4_LUT_B_values_12_port, 
      Inst_clb_slice_4xLUT4_LUT_B_values_13_port, 
      Inst_clb_slice_4xLUT4_LUT_B_values_14_port, 
      Inst_clb_slice_4xLUT4_LUT_B_values_15_port, 
      Inst_clb_slice_4xLUT4_LUT_A_values_0_port, 
      Inst_clb_slice_4xLUT4_LUT_A_values_1_port, 
      Inst_clb_slice_4xLUT4_LUT_A_values_2_port, 
      Inst_clb_slice_4xLUT4_LUT_A_values_3_port, 
      Inst_clb_slice_4xLUT4_LUT_A_values_4_port, 
      Inst_clb_slice_4xLUT4_LUT_A_values_5_port, 
      Inst_clb_slice_4xLUT4_LUT_A_values_6_port, 
      Inst_clb_slice_4xLUT4_LUT_A_values_7_port, 
      Inst_clb_slice_4xLUT4_LUT_A_values_8_port, 
      Inst_clb_slice_4xLUT4_LUT_A_values_9_port, 
      Inst_clb_slice_4xLUT4_LUT_A_values_10_port, 
      Inst_clb_slice_4xLUT4_LUT_A_values_11_port, 
      Inst_clb_slice_4xLUT4_LUT_A_values_12_port, 
      Inst_clb_slice_4xLUT4_LUT_A_values_13_port, 
      Inst_clb_slice_4xLUT4_LUT_A_values_14_port, 
      Inst_clb_slice_4xLUT4_LUT_A_values_15_port, 
      Inst_CLB_switch_matrix_ConfigBits_0_port, 
      Inst_CLB_switch_matrix_ConfigBits_1_port, 
      Inst_CLB_switch_matrix_ConfigBits_2_port, 
      Inst_CLB_switch_matrix_ConfigBits_3_port, 
      Inst_CLB_switch_matrix_ConfigBits_4_port, 
      Inst_CLB_switch_matrix_ConfigBits_5_port, 
      Inst_CLB_switch_matrix_ConfigBits_6_port, 
      Inst_CLB_switch_matrix_ConfigBits_7_port, 
      Inst_CLB_switch_matrix_ConfigBits_8_port, 
      Inst_CLB_switch_matrix_ConfigBits_9_port, 
      Inst_CLB_switch_matrix_ConfigBits_10_port, 
      Inst_CLB_switch_matrix_ConfigBits_11_port, 
      Inst_CLB_switch_matrix_ConfigBits_12_port, 
      Inst_CLB_switch_matrix_ConfigBits_13_port, 
      Inst_CLB_switch_matrix_ConfigBits_14_port, 
      Inst_CLB_switch_matrix_ConfigBits_15_port, 
      Inst_CLB_switch_matrix_ConfigBits_16_port, 
      Inst_CLB_switch_matrix_ConfigBits_17_port, 
      Inst_CLB_switch_matrix_ConfigBits_18_port, 
      Inst_CLB_switch_matrix_ConfigBits_19_port, 
      Inst_CLB_switch_matrix_ConfigBits_20_port, 
      Inst_CLB_switch_matrix_ConfigBits_21_port, 
      Inst_CLB_switch_matrix_ConfigBits_22_port, 
      Inst_CLB_switch_matrix_ConfigBits_23_port, 
      Inst_CLB_switch_matrix_ConfigBits_24_port, 
      Inst_CLB_switch_matrix_ConfigBits_25_port, 
      Inst_CLB_switch_matrix_ConfigBits_26_port, 
      Inst_CLB_switch_matrix_ConfigBits_27_port, 
      Inst_CLB_switch_matrix_ConfigBits_28_port, 
      Inst_CLB_switch_matrix_ConfigBits_29_port, 
      Inst_CLB_switch_matrix_ConfigBits_30_port, 
      Inst_CLB_switch_matrix_ConfigBits_31_port, 
      Inst_CLB_switch_matrix_ConfigBits_32_port, 
      Inst_CLB_switch_matrix_ConfigBits_33_port, 
      Inst_CLB_switch_matrix_ConfigBits_34_port, 
      Inst_CLB_switch_matrix_ConfigBits_35_port, 
      Inst_CLB_switch_matrix_ConfigBits_36_port, 
      Inst_CLB_switch_matrix_ConfigBits_37_port, 
      Inst_CLB_switch_matrix_ConfigBits_38_port, 
      Inst_CLB_switch_matrix_ConfigBits_39_port, 
      Inst_CLB_switch_matrix_ConfigBits_40_port, 
      Inst_CLB_switch_matrix_ConfigBits_41_port, 
      Inst_CLB_switch_matrix_ConfigBits_42_port, 
      Inst_CLB_switch_matrix_ConfigBits_43_port, 
      Inst_CLB_switch_matrix_ConfigBits_44_port, 
      Inst_CLB_switch_matrix_ConfigBits_45_port, 
      Inst_CLB_switch_matrix_ConfigBits_46_port, 
      Inst_CLB_switch_matrix_ConfigBits_47_port, 
      Inst_CLB_switch_matrix_ConfigBits_48_port, 
      Inst_CLB_switch_matrix_ConfigBits_49_port, 
      Inst_CLB_switch_matrix_ConfigBits_50_port, 
      Inst_CLB_switch_matrix_ConfigBits_51_port, 
      Inst_CLB_switch_matrix_ConfigBits_52_port, 
      Inst_CLB_switch_matrix_ConfigBits_53_port, 
      Inst_CLB_switch_matrix_ConfigBits_54_port, 
      Inst_CLB_switch_matrix_ConfigBits_55_port, 
      Inst_CLB_switch_matrix_ConfigBits_56_port, 
      Inst_CLB_switch_matrix_ConfigBits_57_port, 
      Inst_CLB_switch_matrix_ConfigBits_58_port, 
      Inst_CLB_switch_matrix_ConfigBits_59_port, 
      Inst_CLB_switch_matrix_ConfigBits_60_port, 
      Inst_CLB_switch_matrix_ConfigBits_61_port, 
      Inst_CLB_switch_matrix_ConfigBits_62_port, 
      Inst_CLB_switch_matrix_ConfigBits_63_port, 
      Inst_CLB_switch_matrix_ConfigBits_64_port, 
      Inst_CLB_switch_matrix_ConfigBits_65_port, 
      Inst_CLB_switch_matrix_ConfigBits_66_port, 
      Inst_CLB_switch_matrix_ConfigBits_67_port, 
      Inst_CLB_switch_matrix_ConfigBits_68_port, 
      Inst_CLB_switch_matrix_ConfigBits_69_port, 
      Inst_CLB_switch_matrix_ConfigBits_70_port, 
      Inst_CLB_switch_matrix_ConfigBits_71_port, 
      Inst_CLB_switch_matrix_ConfigBits_72_port, 
      Inst_CLB_switch_matrix_ConfigBits_73_port, 
      Inst_CLB_switch_matrix_ConfigBits_74_port, 
      Inst_CLB_switch_matrix_ConfigBits_75_port, 
      Inst_CLB_switch_matrix_ConfigBits_76_port, 
      Inst_CLB_switch_matrix_ConfigBits_77_port, 
      Inst_CLB_switch_matrix_ConfigBits_78_port, 
      Inst_CLB_switch_matrix_ConfigBits_79_port, 
      Inst_CLB_switch_matrix_ConfigBits_80_port, 
      Inst_CLB_switch_matrix_ConfigBits_81_port, 
      Inst_CLB_switch_matrix_ConfigBits_82_port, 
      Inst_CLB_switch_matrix_ConfigBits_83_port, 
      Inst_CLB_switch_matrix_ConfigBits_84_port, 
      Inst_CLB_switch_matrix_ConfigBits_85_port, 
      Inst_CLB_switch_matrix_ConfigBits_86_port, 
      Inst_CLB_switch_matrix_ConfigBits_87_port, 
      Inst_CLB_switch_matrix_ConfigBits_88_port, 
      Inst_CLB_switch_matrix_ConfigBits_89_port, 
      Inst_CLB_switch_matrix_ConfigBits_90_port, 
      Inst_CLB_switch_matrix_ConfigBits_91_port, 
      Inst_CLB_switch_matrix_ConfigBits_92_port, 
      Inst_CLB_switch_matrix_ConfigBits_93_port, 
      Inst_CLB_switch_matrix_ConfigBits_94_port, 
      Inst_CLB_switch_matrix_ConfigBits_95_port, 
      Inst_CLB_switch_matrix_ConfigBits_96_port, 
      Inst_CLB_switch_matrix_ConfigBits_97_port, 
      Inst_CLB_switch_matrix_ConfigBits_98_port, 
      Inst_CLB_switch_matrix_ConfigBits_99_port, 
      Inst_CLB_switch_matrix_ConfigBits_100_port, 
      Inst_CLB_switch_matrix_ConfigBits_101_port, 
      Inst_CLB_switch_matrix_ConfigBits_102_port, 
      Inst_CLB_switch_matrix_ConfigBits_103_port, 
      Inst_CLB_switch_matrix_ConfigBits_104_port, 
      Inst_CLB_switch_matrix_ConfigBits_105_port, 
      Inst_CLB_switch_matrix_ConfigBits_106_port, 
      Inst_CLB_switch_matrix_ConfigBits_107_port, 
      Inst_CLB_switch_matrix_ConfigBits_108_port, 
      Inst_CLB_switch_matrix_ConfigBits_109_port, 
      Inst_CLB_switch_matrix_ConfigBits_110_port, 
      Inst_CLB_switch_matrix_ConfigBits_111_port, 
      Inst_CLB_switch_matrix_ConfigBits_112_port, 
      Inst_CLB_switch_matrix_ConfigBits_113_port, 
      Inst_CLB_switch_matrix_ConfigBits_114_port, 
      Inst_CLB_switch_matrix_ConfigBits_115_port, 
      Inst_CLB_switch_matrix_ConfigBits_116_port, 
      Inst_CLB_switch_matrix_ConfigBits_117_port, 
      Inst_CLB_switch_matrix_ConfigBits_118_port, 
      Inst_CLB_switch_matrix_ConfigBits_119_port, 
      Inst_CLB_switch_matrix_ConfigBits_120_port, 
      Inst_CLB_switch_matrix_ConfigBits_121_port, 
      Inst_CLB_switch_matrix_ConfigBits_122_port, 
      Inst_CLB_switch_matrix_ConfigBits_123_port, 
      Inst_CLB_switch_matrix_ConfigBits_124_port, 
      Inst_CLB_switch_matrix_ConfigBits_125_port, 
      Inst_CLB_switch_matrix_ConfigBits_126_port, 
      Inst_CLB_switch_matrix_ConfigBits_127_port, 
      Inst_CLB_switch_matrix_ConfigBits_128_port, 
      Inst_CLB_switch_matrix_ConfigBits_129_port, 
      Inst_CLB_switch_matrix_ConfigBits_130_port, 
      Inst_CLB_switch_matrix_ConfigBits_131_port, 
      Inst_CLB_switch_matrix_ConfigBits_132_port, 
      Inst_CLB_switch_matrix_ConfigBits_133_port, 
      Inst_CLB_switch_matrix_ConfigBits_134_port, 
      Inst_CLB_switch_matrix_ConfigBits_135_port, 
      Inst_CLB_switch_matrix_ConfigBits_136_port, 
      Inst_CLB_switch_matrix_ConfigBits_137_port, 
      Inst_CLB_switch_matrix_ConfigBits_138_port, 
      Inst_CLB_switch_matrix_ConfigBits_139_port, 
      Inst_CLB_switch_matrix_ConfigBits_140_port, 
      Inst_CLB_switch_matrix_ConfigBits_141_port, 
      Inst_CLB_switch_matrix_ConfigBits_142_port, 
      Inst_CLB_switch_matrix_ConfigBits_143_port, 
      Inst_CLB_switch_matrix_ConfigBits_144_port, 
      Inst_CLB_switch_matrix_ConfigBits_145_port, 
      Inst_CLB_switch_matrix_ConfigBits_146_port, 
      Inst_CLB_switch_matrix_ConfigBits_147_port, 
      Inst_CLB_switch_matrix_ConfigBits_148_port, 
      Inst_CLB_switch_matrix_ConfigBits_149_port, 
      Inst_CLB_switch_matrix_ConfigBits_150_port, 
      Inst_CLB_switch_matrix_ConfigBits_151_port, 
      Inst_CLB_switch_matrix_ConfigBits_152_port, 
      Inst_CLB_switch_matrix_ConfigBits_153_port, 
      Inst_CLB_switch_matrix_ConfigBits_154_port, 
      Inst_CLB_switch_matrix_ConfigBits_155_port, 
      Inst_CLB_switch_matrix_ConfigBits_156_port, 
      Inst_CLB_switch_matrix_ConfigBits_157_port, 
      Inst_CLB_switch_matrix_ConfigBits_158_port, 
      Inst_CLB_switch_matrix_ConfigBits_159_port, 
      Inst_CLB_switch_matrix_ConfigBits_160_port, 
      Inst_CLB_switch_matrix_ConfigBits_161_port, 
      Inst_CLB_switch_matrix_ConfigBits_162_port, 
      Inst_CLB_switch_matrix_ConfigBits_163_port, 
      Inst_CLB_switch_matrix_ConfigBits_164_port, 
      Inst_CLB_switch_matrix_ConfigBits_165_port, 
      Inst_CLB_switch_matrix_ConfigBits_166_port, 
      Inst_CLB_switch_matrix_ConfigBits_167_port, 
      Inst_CLB_switch_matrix_ConfigBits_168_port, 
      Inst_CLB_switch_matrix_ConfigBits_169_port, 
      Inst_CLB_switch_matrix_ConfigBits_170_port, 
      Inst_CLB_switch_matrix_ConfigBits_171_port, 
      Inst_CLB_switch_matrix_ConfigBits_172_port, 
      Inst_CLB_switch_matrix_ConfigBits_173_port, 
      Inst_CLB_switch_matrix_ConfigBits_174_port, 
      Inst_CLB_switch_matrix_ConfigBits_175_port, 
      Inst_CLB_switch_matrix_ConfigBits_176_port, 
      Inst_CLB_switch_matrix_ConfigBits_177_port, 
      Inst_CLB_switch_matrix_ConfigBits_178_port, 
      Inst_CLB_switch_matrix_ConfigBits_179_port, 
      Inst_CLB_switch_matrix_ConfigBits_180_port, n118, n121, n123, n126, n127,
      n129, n130, n134, n135, n136, n137, n138, n140, n203, n218, n270, n464, 
      n505, n506, n507, n509, n513, n514, n515, n516, n517, n518, n520, n521, 
      n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, 
      n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, 
      n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, 
      n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, 
      n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, 
      n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, 
      n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, 
      n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, 
      n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, 
      n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, 
      n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, 
      n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, 
      n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, 
      n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, 
      n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, 
      n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, 
      n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, 
      n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, 
      n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, 
      n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, 
      n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, 
      n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, 
      n795, n797, n799, n800, n801, n802, n804, n805, n806, n807, n808, n810, 
      n812, n814, n816, n818, n820, n822, n824, n826, n828, n830, n832, n834, 
      n836, n838, n840, n842, n844, n846, n848, n850, n852, n854, n856, n857, 
      n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, 
      n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, 
      n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, 
      n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, 
      n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, 
      n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, 
      n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, 
      n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, 
      n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, 
      n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, 
      n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, 
      n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002
      , n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, 
      n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, 
      n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, 
      n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, 
      n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, 
      n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, 
      n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, 
      n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, 
      n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, 
      n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, 
      n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, 
      n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, 
      n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, 
      n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, 
      n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, 
      n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, 
      n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, 
      n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, 
      n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, 
      n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, 
      n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, 
      n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, 
      n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, 
      n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, 
      n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, 
      n1253, n1254, n1255, n1256, n1257 : std_logic;

begin
   
   Inst_test_C17 : XOR2D1 port map( A1 => TestIn, A2 => conf_data_2_port, Z => 
                           TestOut);
   Inst_clb_slice_4xLUT4_LUT_A_values_reg_0_inst : DFQD1 port map( D => n776, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_A_values_0_port);
   Inst_clb_slice_4xLUT4_LUT_A_values_reg_1_inst : DFQD1 port map( D => n775, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_A_values_1_port);
   Inst_clb_slice_4xLUT4_LUT_A_values_reg_2_inst : DFQD1 port map( D => n774, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_A_values_2_port);
   Inst_clb_slice_4xLUT4_LUT_A_values_reg_3_inst : DFQD1 port map( D => n773, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_A_values_3_port);
   Inst_clb_slice_4xLUT4_LUT_A_values_reg_4_inst : DFQD1 port map( D => n772, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_A_values_4_port);
   Inst_clb_slice_4xLUT4_LUT_A_values_reg_5_inst : DFQD1 port map( D => n771, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_A_values_5_port);
   Inst_clb_slice_4xLUT4_LUT_A_values_reg_6_inst : DFQD1 port map( D => n770, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_A_values_6_port);
   Inst_clb_slice_4xLUT4_LUT_A_values_reg_7_inst : DFQD1 port map( D => n769, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_A_values_7_port);
   Inst_clb_slice_4xLUT4_LUT_A_values_reg_8_inst : DFQD1 port map( D => n768, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_A_values_8_port);
   Inst_clb_slice_4xLUT4_LUT_A_values_reg_9_inst : DFQD1 port map( D => n767, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_A_values_9_port);
   Inst_clb_slice_4xLUT4_LUT_A_values_reg_10_inst : DFQD1 port map( D => n766, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_A_values_10_port);
   Inst_clb_slice_4xLUT4_LUT_A_values_reg_11_inst : DFQD1 port map( D => n765, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_A_values_11_port);
   Inst_clb_slice_4xLUT4_LUT_A_values_reg_12_inst : DFQD1 port map( D => n764, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_A_values_12_port);
   Inst_clb_slice_4xLUT4_LUT_A_values_reg_13_inst : DFQD1 port map( D => n763, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_A_values_13_port);
   Inst_clb_slice_4xLUT4_LUT_A_values_reg_14_inst : DFQD1 port map( D => n762, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_A_values_14_port);
   Inst_clb_slice_4xLUT4_LUT_A_values_reg_15_inst : DFQD1 port map( D => n761, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_A_values_15_port);
   Inst_clb_slice_4xLUT4_LUT_B_values_reg_0_inst : DFQD1 port map( D => n760, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_B_values_0_port);
   Inst_clb_slice_4xLUT4_LUT_B_values_reg_1_inst : DFQD1 port map( D => n759, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_B_values_1_port);
   Inst_clb_slice_4xLUT4_LUT_B_values_reg_2_inst : DFQD1 port map( D => n758, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_B_values_2_port);
   Inst_clb_slice_4xLUT4_LUT_B_values_reg_3_inst : DFQD1 port map( D => n757, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_B_values_3_port);
   Inst_clb_slice_4xLUT4_LUT_B_values_reg_4_inst : DFQD1 port map( D => n756, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_B_values_4_port);
   Inst_clb_slice_4xLUT4_LUT_B_values_reg_5_inst : DFQD1 port map( D => n755, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_B_values_5_port);
   Inst_clb_slice_4xLUT4_LUT_B_values_reg_6_inst : DFQD1 port map( D => n754, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_B_values_6_port);
   Inst_clb_slice_4xLUT4_LUT_B_values_reg_7_inst : DFQD1 port map( D => n753, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_B_values_7_port);
   Inst_clb_slice_4xLUT4_LUT_B_values_reg_8_inst : DFQD1 port map( D => n752, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_B_values_8_port);
   Inst_clb_slice_4xLUT4_LUT_B_values_reg_9_inst : DFQD1 port map( D => n751, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_B_values_9_port);
   Inst_clb_slice_4xLUT4_LUT_B_values_reg_10_inst : DFQD1 port map( D => n750, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_B_values_10_port);
   Inst_clb_slice_4xLUT4_LUT_B_values_reg_11_inst : DFQD1 port map( D => n749, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_B_values_11_port);
   Inst_clb_slice_4xLUT4_LUT_B_values_reg_12_inst : DFQD1 port map( D => n748, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_B_values_12_port);
   Inst_clb_slice_4xLUT4_LUT_B_values_reg_13_inst : DFQD1 port map( D => n747, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_B_values_13_port);
   Inst_clb_slice_4xLUT4_LUT_B_values_reg_14_inst : DFQD1 port map( D => n746, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_B_values_14_port);
   Inst_clb_slice_4xLUT4_LUT_B_values_reg_15_inst : DFQD1 port map( D => n745, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_B_values_15_port);
   Inst_clb_slice_4xLUT4_LUT_C_values_reg_0_inst : DFQD1 port map( D => n744, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_C_values_0_port);
   Inst_clb_slice_4xLUT4_LUT_C_values_reg_1_inst : DFQD1 port map( D => n743, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_C_values_1_port);
   Inst_clb_slice_4xLUT4_LUT_C_values_reg_2_inst : DFQD1 port map( D => n742, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_C_values_2_port);
   Inst_clb_slice_4xLUT4_LUT_C_values_reg_3_inst : DFQD1 port map( D => n741, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_C_values_3_port);
   Inst_clb_slice_4xLUT4_LUT_C_values_reg_4_inst : DFQD1 port map( D => n740, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_C_values_4_port);
   Inst_clb_slice_4xLUT4_LUT_C_values_reg_5_inst : DFQD1 port map( D => n739, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_C_values_5_port);
   Inst_clb_slice_4xLUT4_LUT_C_values_reg_6_inst : DFQD1 port map( D => n738, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_C_values_6_port);
   Inst_clb_slice_4xLUT4_LUT_C_values_reg_7_inst : DFQD1 port map( D => n737, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_C_values_7_port);
   Inst_clb_slice_4xLUT4_LUT_C_values_reg_8_inst : DFQD1 port map( D => n736, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_C_values_8_port);
   Inst_clb_slice_4xLUT4_LUT_C_values_reg_9_inst : DFQD1 port map( D => n735, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_C_values_9_port);
   Inst_clb_slice_4xLUT4_LUT_C_values_reg_10_inst : DFQD1 port map( D => n734, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_C_values_10_port);
   Inst_clb_slice_4xLUT4_LUT_C_values_reg_11_inst : DFQD1 port map( D => n733, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_C_values_11_port);
   Inst_clb_slice_4xLUT4_LUT_C_values_reg_12_inst : DFQD1 port map( D => n732, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_C_values_12_port);
   Inst_clb_slice_4xLUT4_LUT_C_values_reg_13_inst : DFQD1 port map( D => n731, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_C_values_13_port);
   Inst_clb_slice_4xLUT4_LUT_C_values_reg_14_inst : DFQD1 port map( D => n730, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_C_values_14_port);
   Inst_clb_slice_4xLUT4_LUT_C_values_reg_15_inst : DFQD1 port map( D => n729, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_C_values_15_port);
   Inst_clb_slice_4xLUT4_LUT_D_values_reg_0_inst : DFQD1 port map( D => n728, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_D_values_0_port);
   Inst_clb_slice_4xLUT4_LUT_D_values_reg_1_inst : DFQD1 port map( D => n727, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_D_values_1_port);
   Inst_clb_slice_4xLUT4_LUT_D_values_reg_2_inst : DFQD1 port map( D => n726, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_D_values_2_port);
   Inst_clb_slice_4xLUT4_LUT_D_values_reg_3_inst : DFQD1 port map( D => n725, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_D_values_3_port);
   Inst_clb_slice_4xLUT4_LUT_D_values_reg_4_inst : DFQD1 port map( D => n724, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_D_values_4_port);
   Inst_clb_slice_4xLUT4_LUT_D_values_reg_5_inst : DFQD1 port map( D => n723, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_D_values_5_port);
   Inst_clb_slice_4xLUT4_LUT_D_values_reg_6_inst : DFQD1 port map( D => n722, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_D_values_6_port);
   Inst_clb_slice_4xLUT4_LUT_D_values_reg_7_inst : DFQD1 port map( D => n721, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_D_values_7_port);
   Inst_clb_slice_4xLUT4_LUT_D_values_reg_8_inst : DFQD1 port map( D => n720, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_D_values_8_port);
   Inst_clb_slice_4xLUT4_LUT_D_values_reg_9_inst : DFQD1 port map( D => n719, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_D_values_9_port);
   Inst_clb_slice_4xLUT4_LUT_D_values_reg_10_inst : DFQD1 port map( D => n718, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_D_values_10_port);
   Inst_clb_slice_4xLUT4_LUT_D_values_reg_11_inst : DFQD1 port map( D => n717, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_D_values_11_port);
   Inst_clb_slice_4xLUT4_LUT_D_values_reg_12_inst : DFQD1 port map( D => n716, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_D_values_12_port);
   Inst_clb_slice_4xLUT4_LUT_D_values_reg_13_inst : DFQD1 port map( D => n715, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_D_values_13_port);
   Inst_clb_slice_4xLUT4_LUT_D_values_reg_14_inst : DFQD1 port map( D => n714, 
                           CP => CLK, Q => 
                           Inst_clb_slice_4xLUT4_LUT_D_values_14_port);
   Inst_clb_slice_4xLUT4_LUT_D_values_reg_15_inst : DFQD1 port map( D => n713, 
                           CP => CLK, Q => conf_data_1_port);
   Inst_test_congig_bit_reg : DFQD1 port map( D => n712, CP => CLK, Q => 
                           conf_data_2_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_180_inst : DFQD1 port map( D => n710, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_180_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_179_inst : DFQD1 port map( D => n709, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_179_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_178_inst : DFQD1 port map( D => n708, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_178_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_177_inst : DFQD1 port map( D => n707, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_177_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_176_inst : DFQD1 port map( D => n706, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_176_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_175_inst : DFQD1 port map( D => n705, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_175_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_172_inst : DFQD1 port map( D => n702, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_172_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_170_inst : DFQD1 port map( D => n700, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_170_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_169_inst : DFQD1 port map( D => n699, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_169_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_168_inst : DFQD1 port map( D => n698, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_168_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_167_inst : DFQD1 port map( D => n697, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_167_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_166_inst : DFQD1 port map( D => n696, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_166_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_165_inst : DFQD1 port map( D => n695, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_165_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_164_inst : DFQD1 port map( D => n694, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_164_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_163_inst : DFQD1 port map( D => n693, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_163_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_162_inst : DFQD1 port map( D => n692, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_162_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_160_inst : DFQD1 port map( D => n690, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_160_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_158_inst : DFQD1 port map( D => n688, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_158_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_157_inst : DFQD1 port map( D => n687, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_157_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_155_inst : DFQD1 port map( D => n685, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_155_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_154_inst : DFQD1 port map( D => n684, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_154_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_152_inst : DFQD1 port map( D => n682, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_152_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_151_inst : DFQD1 port map( D => n681, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_151_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_150_inst : DFQD1 port map( D => n680, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_150_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_149_inst : DFQD1 port map( D => n679, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_149_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_147_inst : DFQD1 port map( D => n677, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_147_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_146_inst : DFQD1 port map( D => n676, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_146_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_145_inst : DFQD1 port map( D => n675, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_145_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_143_inst : DFQD1 port map( D => n673, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_143_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_141_inst : DFQD1 port map( D => n671, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_141_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_139_inst : DFQD1 port map( D => n669, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_139_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_137_inst : DFQD1 port map( D => n667, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_137_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_136_inst : DFQD1 port map( D => n666, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_136_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_135_inst : DFQD1 port map( D => n665, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_135_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_134_inst : DFQD1 port map( D => n664, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_134_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_133_inst : DFQD1 port map( D => n663, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_133_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_132_inst : DFQD1 port map( D => n662, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_132_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_131_inst : DFQD1 port map( D => n661, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_131_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_130_inst : DFQD1 port map( D => n660, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_130_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_129_inst : DFQD1 port map( D => n659, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_129_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_128_inst : DFQD1 port map( D => n658, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_128_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_127_inst : DFQD1 port map( D => n657, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_127_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_126_inst : DFQD1 port map( D => n656, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_126_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_125_inst : DFQD1 port map( D => n655, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_125_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_124_inst : DFQD1 port map( D => n654, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_124_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_123_inst : DFQD1 port map( D => n653, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_123_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_122_inst : DFQD1 port map( D => n652, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_122_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_121_inst : DFQD1 port map( D => n651, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_121_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_120_inst : DFQD1 port map( D => n650, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_120_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_119_inst : DFQD1 port map( D => n649, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_119_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_118_inst : DFQD1 port map( D => n648, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_118_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_117_inst : DFQD1 port map( D => n647, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_117_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_116_inst : DFQD1 port map( D => n646, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_116_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_115_inst : DFQD1 port map( D => n645, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_115_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_113_inst : DFQD1 port map( D => n643, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_113_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_112_inst : DFQD1 port map( D => n642, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_112_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_111_inst : DFQD1 port map( D => n641, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_111_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_110_inst : DFQD1 port map( D => n640, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_110_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_109_inst : DFQD1 port map( D => n639, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_109_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_108_inst : DFQD1 port map( D => n638, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_108_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_107_inst : DFQD1 port map( D => n637, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_107_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_106_inst : DFQD1 port map( D => n636, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_106_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_105_inst : DFQD1 port map( D => n635, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_105_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_104_inst : DFQD1 port map( D => n634, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_104_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_103_inst : DFQD1 port map( D => n633, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_103_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_102_inst : DFQD1 port map( D => n632, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_102_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_101_inst : DFQD1 port map( D => n631, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_101_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_100_inst : DFQD1 port map( D => n630, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_100_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_99_inst : DFQD1 port map( D => n629, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_99_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_98_inst : DFQD1 port map( D => n628, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_98_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_97_inst : DFQD1 port map( D => n627, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_97_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_96_inst : DFQD1 port map( D => n626, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_96_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_95_inst : DFQD1 port map( D => n625, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_95_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_94_inst : DFQD1 port map( D => n624, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_94_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_93_inst : DFQD1 port map( D => n623, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_93_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_92_inst : DFQD1 port map( D => n622, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_92_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_91_inst : DFQD1 port map( D => n621, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_91_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_90_inst : DFQD1 port map( D => n620, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_90_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_89_inst : DFQD1 port map( D => n619, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_89_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_88_inst : DFQD1 port map( D => n618, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_88_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_87_inst : DFQD1 port map( D => n617, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_87_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_86_inst : DFQD1 port map( D => n616, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_86_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_85_inst : DFQD1 port map( D => n615, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_85_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_84_inst : DFQD1 port map( D => n614, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_84_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_83_inst : DFQD1 port map( D => n613, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_83_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_82_inst : DFQD1 port map( D => n612, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_82_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_81_inst : DFQD1 port map( D => n611, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_81_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_80_inst : DFQD1 port map( D => n610, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_80_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_79_inst : DFQD1 port map( D => n609, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_79_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_78_inst : DFQD1 port map( D => n608, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_78_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_77_inst : DFQD1 port map( D => n607, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_77_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_76_inst : DFQD1 port map( D => n606, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_76_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_75_inst : DFQD1 port map( D => n605, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_75_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_74_inst : DFQD1 port map( D => n604, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_74_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_73_inst : DFQD1 port map( D => n603, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_73_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_72_inst : DFQD1 port map( D => n602, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_72_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_71_inst : DFQD1 port map( D => n601, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_71_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_70_inst : DFQD1 port map( D => n600, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_70_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_69_inst : DFQD1 port map( D => n599, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_69_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_68_inst : DFQD1 port map( D => n598, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_68_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_67_inst : DFQD1 port map( D => n597, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_67_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_66_inst : DFQD1 port map( D => n596, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_66_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_65_inst : DFQD1 port map( D => n595, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_65_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_64_inst : DFQD1 port map( D => n594, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_64_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_63_inst : DFQD1 port map( D => n593, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_63_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_62_inst : DFQD1 port map( D => n592, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_62_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_61_inst : DFQD1 port map( D => n591, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_61_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_60_inst : DFQD1 port map( D => n590, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_60_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_59_inst : DFQD1 port map( D => n589, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_59_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_58_inst : DFQD1 port map( D => n588, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_58_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_57_inst : DFQD1 port map( D => n587, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_57_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_56_inst : DFQD1 port map( D => n586, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_56_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_55_inst : DFQD1 port map( D => n585, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_55_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_54_inst : DFQD1 port map( D => n584, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_54_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_53_inst : DFQD1 port map( D => n583, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_53_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_52_inst : DFQD1 port map( D => n582, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_52_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_51_inst : DFQD1 port map( D => n581, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_51_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_50_inst : DFQD1 port map( D => n580, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_50_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_49_inst : DFQD1 port map( D => n579, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_49_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_48_inst : DFQD1 port map( D => n578, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_48_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_47_inst : DFQD1 port map( D => n577, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_47_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_46_inst : DFQD1 port map( D => n576, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_46_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_45_inst : DFQD1 port map( D => n575, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_45_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_44_inst : DFQD1 port map( D => n574, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_44_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_43_inst : DFQD1 port map( D => n573, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_43_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_42_inst : DFQD1 port map( D => n572, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_42_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_41_inst : DFQD1 port map( D => n571, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_41_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_40_inst : DFQD1 port map( D => n570, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_40_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_39_inst : DFQD1 port map( D => n569, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_39_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_38_inst : DFQD1 port map( D => n568, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_38_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_37_inst : DFQD1 port map( D => n567, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_37_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_36_inst : DFQD1 port map( D => n566, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_36_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_35_inst : DFQD1 port map( D => n565, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_35_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_34_inst : DFQD1 port map( D => n564, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_34_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_33_inst : DFQD1 port map( D => n563, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_33_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_32_inst : DFQD1 port map( D => n562, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_32_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_31_inst : DFQD1 port map( D => n561, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_31_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_30_inst : DFQD1 port map( D => n560, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_30_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_29_inst : DFQD1 port map( D => n559, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_29_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_28_inst : DFQD1 port map( D => n558, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_28_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_27_inst : DFQD1 port map( D => n557, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_27_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_26_inst : DFQD1 port map( D => n556, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_26_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_25_inst : DFQD1 port map( D => n555, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_25_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_24_inst : DFQD1 port map( D => n554, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_24_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_23_inst : DFQD1 port map( D => n553, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_23_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_22_inst : DFQD1 port map( D => n552, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_22_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_21_inst : DFQD1 port map( D => n551, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_21_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_20_inst : DFQD1 port map( D => n550, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_20_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_19_inst : DFQD1 port map( D => n549, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_19_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_18_inst : DFQD1 port map( D => n548, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_18_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_17_inst : DFQD1 port map( D => n547, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_17_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_16_inst : DFQD1 port map( D => n546, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_16_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_15_inst : DFQD1 port map( D => n545, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_15_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_14_inst : DFQD1 port map( D => n544, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_14_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_13_inst : DFQD1 port map( D => n543, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_13_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_12_inst : DFQD1 port map( D => n542, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_12_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_11_inst : DFQD1 port map( D => n541, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_11_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_10_inst : DFQD1 port map( D => n540, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_10_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_9_inst : DFQD1 port map( D => n539, CP
                           => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_9_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_8_inst : DFQD1 port map( D => n538, CP
                           => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_8_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_7_inst : DFQD1 port map( D => n537, CP
                           => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_7_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_6_inst : DFQD1 port map( D => n536, CP
                           => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_6_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_5_inst : DFQD1 port map( D => n535, CP
                           => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_5_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_4_inst : DFQD1 port map( D => n534, CP
                           => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_4_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_3_inst : DFQD1 port map( D => n533, CP
                           => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_3_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_2_inst : DFQD1 port map( D => n532, CP
                           => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_2_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_1_inst : DFQD1 port map( D => n531, CP
                           => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_1_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_0_inst : DFQD1 port map( D => n530, CP
                           => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_0_port);
   U497 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_177_port, 
                           A2 => n270, B1 => n515, B2 => n118, ZN => 
                           IJ_BEG_11_port);
   U502 : AOI22D1 port map( A1 => n857, A2 => n218, B1 => n529, B2 => n856, ZN 
                           => OJ_BEG_2_port);
   U504 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_153_port, 
                           A2 => IJ_BEG_11_port, B1 => D, B2 => n121, ZN => 
                           n123);
   U509 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_171_port, 
                           A2 => n514, B1 => n518, B2 => n127, ZN => n126);
   U511 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_171_port, 
                           A2 => n218, B1 => n203, B2 => n127, ZN => n130);
   U514 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_171_port, 
                           A2 => n517, B1 => n464, B2 => n127, ZN => n129);
   U518 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_159_port, 
                           A2 => OJ_BEG_0_port, B1 => TestOut, B2 => n135, ZN 
                           => n134);
   U519 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_161_port, 
                           A2 => n526, B1 => n134, B2 => n136, ZN => n140);
   U520 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_159_port, 
                           A2 => OJ_BEG_2_port, B1 => OJ_BEG_1_port, B2 => n135
                           , ZN => n138);
   U521 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_159_port, 
                           A2 => DQ, B1 => D, B2 => n135, ZN => n137);
   U819 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_156_port, 
                           A2 => OJ_BEG_2_port, B1 => OJ_BEG_1_port, B2 => n505
                           , ZN => n513);
   U821 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_156_port, 
                           A2 => n507, B1 => n506, B2 => n505, ZN => n509);
   U824 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_174_port, 
                           A2 => n515, B1 => n514, B2 => n516, ZN => n521);
   U825 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_174_port, 
                           A2 => n518, B1 => n517, B2 => n516, ZN => n520);
   U827 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_176_port, 
                           A2 => n525, B1 => n523, B2 => n522, ZN => 
                           IJ_BEG_10_port);
   U828 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_179_port, 
                           A2 => n526, B1 => n525, B2 => n524, ZN => 
                           OJ_BEG_0_port);
   U829 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_178_port, 
                           A2 => n529, B1 => n528, B2 => n527, ZN => 
                           IJ_BEG_12_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_114_inst : DFQD1 port map( D => n644, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_114_port);
   Inst_clb_slice_4xLUT4_BQ_reg : DFQD1 port map( D => B, CP => CLK, Q => BQ);
   Inst_clb_slice_4xLUT4_AQ_reg : DFQD1 port map( D => A, CP => CLK, Q => AQ);
   Inst_clb_slice_4xLUT4_CQ_reg : DFQD1 port map( D => C, CP => CLK, Q => CQ);
   Inst_CLB_switch_matrix_ConfigBits_reg_144_inst : DFQD1 port map( D => n674, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_144_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_142_inst : DFQD1 port map( D => n672, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_142_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_140_inst : DFQD1 port map( D => n670, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_140_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_138_inst : DFQD1 port map( D => n668, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_138_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_153_inst : DFQD1 port map( D => n683, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_153_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_148_inst : DFQD1 port map( D => n678, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_148_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_174_inst : DFQD1 port map( D => n704, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_174_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_156_inst : DFQD1 port map( D => n686, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_156_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_171_inst : DFQD1 port map( D => n701, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_171_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_173_inst : DFQD1 port map( D => n703, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_173_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_161_inst : DFQD1 port map( D => n691, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_161_port);
   Inst_clb_slice_4xLUT4_DQ_reg : DFQD1 port map( D => D, CP => CLK, Q => DQ);
   Inst_CLB_switch_matrix_ConfigBits_reg_159_inst : DFQD1 port map( D => n689, 
                           CP => CLK, Q => 
                           Inst_CLB_switch_matrix_ConfigBits_159_port);
   Inst_CLB_switch_matrix_ConfigBits_reg_181_inst : DFQD1 port map( D => n711, 
                           CP => CLK, Q => n1342);
   U830 : MUX4D4 port map( I0 => W2END(3), I1 => W2END(5), I2 => W2END(4), I3 
                           => A, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_108_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_107_port, Z => 
                           n1332);
   U831 : INVD0 port map( I => MODE, ZN => n779);
   U832 : INVD1 port map( I => MODE, ZN => n778);
   U833 : INVD1 port map( I => MODE, ZN => n777);
   U834 : INVD0 port map( I => MODE, ZN => n783);
   U835 : INVD0 port map( I => MODE, ZN => n782);
   U836 : INVD0 port map( I => MODE, ZN => n781);
   U837 : INVD0 port map( I => MODE, ZN => n780);
   U838 : OR2D0 port map( A1 => n954, A2 => n953, Z => n966);
   U839 : OR2D0 port map( A1 => n956, A2 => n955, Z => n965);
   U840 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_116_port, ZN 
                           => n1142);
   U841 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_151_port, ZN 
                           => n1107);
   U842 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_152_port, ZN 
                           => n1106);
   U843 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_154_port, ZN 
                           => n1105);
   U844 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_157_port, ZN 
                           => n1103);
   U845 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_158_port, ZN 
                           => n1102);
   U846 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_165_port, ZN 
                           => n1097);
   U847 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_175_port, ZN 
                           => n1089);
   U848 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_180_port, ZN 
                           => n1088);
   U849 : MUX4ND0 port map( I0 => n985, I1 => n984, I2 => n983, I3 => n982, S0 
                           => Inst_CLB_switch_matrix_ConfigBits_100_port, S1 =>
                           Inst_CLB_switch_matrix_ConfigBits_98_port, ZN => 
                           n1335);
   U850 : INVD0 port map( I => n1334, ZN => n850);
   U851 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_102_port, 
                           A2 => n981, B1 => n980, B2 => n1156, ZN => n1334);
   U852 : INVD0 port map( I => n1333, ZN => n848);
   U853 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_105_port, 
                           A2 => n977, B1 => n976, B2 => n1153, ZN => n1333);
   U854 : INVD0 port map( I => n1331, ZN => n797);
   U855 : INVD0 port map( I => n1330, ZN => n795);
   U856 : INVD0 port map( I => n1329, ZN => n846);
   U857 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_77_port, A2
                           => n1007, B1 => n1006, B2 => n1181, ZN => n1329);
   U858 : INVD0 port map( I => n1328, ZN => n844);
   U859 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_79_port, A2
                           => n1003, B1 => n1002, B2 => n1179, ZN => n1328);
   U860 : MUX4ND0 port map( I0 => n1023, I1 => n1022, I2 => n1021, I3 => n218, 
                           S0 => Inst_CLB_switch_matrix_ConfigBits_88_port, S1 
                           => Inst_CLB_switch_matrix_ConfigBits_86_port, ZN => 
                           n1327);
   U861 : MUX4ND0 port map( I0 => n992, I1 => n991, I2 => n990, I3 => n989, S0 
                           => Inst_CLB_switch_matrix_ConfigBits_92_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_90_port, ZN => 
                           n1326);
   U862 : MUX4ND0 port map( I0 => n900, I1 => n899, I2 => n898, I3 => n897, S0 
                           => Inst_CLB_switch_matrix_ConfigBits_96_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_94_port, ZN => 
                           n1325);
   U863 : INVD0 port map( I => n1319, ZN => n842);
   U864 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_62_port, A2
                           => n998, B1 => n997, B2 => n1196, ZN => n1319);
   U865 : INVD0 port map( I => n1318, ZN => n840);
   U866 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_65_port, A2
                           => n979, B1 => n978, B2 => n1193, ZN => n1318);
   U867 : INVD0 port map( I => n1317, ZN => n838);
   U868 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_68_port, A2
                           => n988, B1 => n987, B2 => n1190, ZN => n1317);
   U869 : MUX4D1 port map( I0 => S2END(3), I1 => S2END(4), I2 => W1END(0), I3 
                           => W1END(1), S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_70_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_71_port, Z => 
                           n1316);
   U870 : INVD0 port map( I => n1315, ZN => n854);
   U871 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_74_port, A2
                           => n270, B1 => n1001, B2 => n1184, ZN => n1315);
   U872 : INVD0 port map( I => n1314, ZN => n836);
   U873 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_47_port, A2
                           => n973, B1 => n972, B2 => n1211, ZN => n1314);
   U874 : INVD0 port map( I => n1313, ZN => n834);
   U875 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_50_port, A2
                           => n969, B1 => n968, B2 => n1208, ZN => n1313);
   U876 : INVD0 port map( I => n1312, ZN => n832);
   U877 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_54_port, A2
                           => n1017, B1 => n1016, B2 => n1204, ZN => n1312);
   U878 : INVD0 port map( I => n1311, ZN => n830);
   U879 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_56_port, A2
                           => n904, B1 => n903, B2 => n1202, ZN => n1311);
   U880 : INVD0 port map( I => n1310, ZN => n828);
   U881 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_59_port, A2
                           => n1013, B1 => n1012, B2 => n1199, ZN => n1310);
   U882 : INVD0 port map( I => n1305, ZN => n852);
   U883 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_36_port, A2
                           => n896, B1 => n895, B2 => n1222, ZN => n1305);
   U884 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_35_port, A2
                           => IJ_BEG_0_port, B1 => n894, B2 => n1223, ZN => 
                           n896);
   U885 : INVD0 port map( I => n1304, ZN => n826);
   U886 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_38_port, A2
                           => n892, B1 => n891, B2 => n1220, ZN => n1304);
   U887 : INVD0 port map( I => n1303, ZN => n824);
   U888 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_41_port, A2
                           => n1005, B1 => n1004, B2 => n1217, ZN => n1303);
   U889 : INVD0 port map( I => n1302, ZN => n822);
   U890 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_44_port, A2
                           => n971, B1 => n970, B2 => n1214, ZN => n1302);
   U891 : INVD0 port map( I => n1301, ZN => n820);
   U892 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_21_port, A2
                           => n890, B1 => n889, B2 => n1237, ZN => n1301);
   U893 : INVD0 port map( I => n1300, ZN => n818);
   U894 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_24_port, A2
                           => n1000, B1 => n999, B2 => n1234, ZN => n1300);
   U895 : AOI221D1 port map( A1 => n887, A2 => 
                           Inst_CLB_switch_matrix_ConfigBits_27_port, B1 => 
                           n886, B2 => n1231, C => 
                           Inst_CLB_switch_matrix_ConfigBits_29_port, ZN => 
                           n888);
   U896 : INVD0 port map( I => n1292, ZN => n816);
   U897 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_16_port, A2
                           => n1020, B1 => n1019, B2 => n1242, ZN => n1292);
   U898 : INVD0 port map( I => n1291, ZN => n814);
   U899 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_18_port, A2
                           => n885, B1 => n884, B2 => n1240, ZN => n1291);
   U900 : MUX4D1 port map( I0 => N2END(0), I1 => N2END(2), I2 => N2END(1), I3 
                           => N4END(0), S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_7_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_6_port, Z => n1287
                           );
   U901 : INVD0 port map( I => n1286, ZN => n812);
   U902 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_10_port, A2
                           => n528, B1 => n986, B2 => n1248, ZN => n1286);
   U903 : INVD0 port map( I => n1285, ZN => n810);
   U904 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_13_port, A2
                           => n975, B1 => n974, B2 => n1245, ZN => n1285);
   U905 : MUX4D1 port map( I0 => N1END(0), I1 => N1END(2), I2 => N1END(1), I3 
                           => N2END(0), S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_1_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_0_port, Z => n1284
                           );
   U906 : MUX4D1 port map( I0 => N1END(1), I1 => N2END(0), I2 => N1END(2), I3 
                           => N2END(1), S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_3_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_2_port, Z => n1283
                           );
   U907 : MUX4D1 port map( I0 => N1END(2), I1 => N2END(1), I2 => N2END(0), I3 
                           => N2END(2), S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_5_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_4_port, Z => n1282
                           );
   U908 : MUX4ND0 port map( I0 => OJ_BEG_1_port, I1 => IJ_BEG_9_port, I2 => 
                           OJ_BEG_2_port, I3 => IJ_BEG_10_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_163_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_162_port, ZN => 
                           n882);
   U909 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_178_port, ZN 
                           => n527);
   U910 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_179_port, ZN 
                           => n524);
   U911 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_176_port, ZN 
                           => n522);
   U912 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_174_port, ZN 
                           => n516);
   U913 : INVD0 port map( I => DQ, ZN => n507);
   U914 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_156_port, ZN 
                           => n505);
   U915 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_161_port, ZN 
                           => n136);
   U916 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_159_port, ZN 
                           => n135);
   U917 : OR2D0 port map( A1 => n870, A2 => n869, Z => n871);
   U918 : OR2D0 port map( A1 => n866, A2 => n865, Z => n872);
   U919 : OR2D0 port map( A1 => n864, A2 => n863, Z => n873);
   U920 : INVD0 port map( I => IJ_BEG_11_port, ZN => n218);
   U921 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_177_port, ZN 
                           => n118);
   U922 : MUX2D0 port map( I0 => Inst_clb_slice_4xLUT4_LUT_A_values_0_port, I1 
                           => CONFin, S => MODE, Z => n776);
   U923 : AO22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_81_port, A2 
                           => n203, B1 => n526, B2 => n1177, Z => n784);
   U924 : AO22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_30_port, A2 
                           => n993, B1 => n218, B2 => n1228, Z => n785);
   U925 : INVD0 port map( I => n1335, ZN => n862);
   U926 : INVD16 port map( I => n862, ZN => W2BEG(6));
   U927 : INVD0 port map( I => n1327, ZN => n861);
   U928 : INVD16 port map( I => n861, ZN => W1BEG(3));
   U929 : INVD0 port map( I => n1326, ZN => n860);
   U930 : INVD16 port map( I => n860, ZN => W1BEG(4));
   U931 : INVD0 port map( I => n1325, ZN => n859);
   U932 : INVD16 port map( I => n859, ZN => W1BEG(5));
   U933 : INVD0 port map( I => n1316, ZN => n808);
   U934 : INVD16 port map( I => n808, ZN => S2BEG(8));
   U935 : INVD0 port map( I => n1284, ZN => n806);
   U936 : INVD16 port map( I => n806, ZN => N1BEG(0));
   U937 : INVD0 port map( I => n1287, ZN => n807);
   U938 : INVD16 port map( I => n807, ZN => N2BEG(3));
   U939 : INVD0 port map( I => n1282, ZN => n804);
   U940 : INVD16 port map( I => n804, ZN => N1BEG(2));
   U941 : INVD0 port map( I => n1283, ZN => n805);
   U942 : INVD16 port map( I => n805, ZN => N1BEG(1));
   U943 : INVD16 port map( I => n795, ZN => W2BEG(11));
   U944 : INVD16 port map( I => n797, ZN => W2BEG(10));
   U945 : INVD16 port map( I => n799, ZN => E1BEG(3));
   U946 : NR2D0 port map( A1 => n785, A2 => n1225, ZN => n800);
   U947 : NR2D1 port map( A1 => n800, A2 => n996, ZN => n799);
   U948 : AOI221D1 port map( A1 => n995, A2 => 
                           Inst_CLB_switch_matrix_ConfigBits_31_port, B1 => 
                           n994, B2 => n1227, C => 
                           Inst_CLB_switch_matrix_ConfigBits_33_port, ZN => 
                           n996);
   U949 : INVD16 port map( I => n801, ZN => W1BEG(2));
   U950 : NR2D0 port map( A1 => n784, A2 => n1174, ZN => n802);
   U951 : NR2D1 port map( A1 => n802, A2 => n1010, ZN => n801);
   U952 : AOI221D1 port map( A1 => n1009, A2 => 
                           Inst_CLB_switch_matrix_ConfigBits_82_port, B1 => 
                           n1008, B2 => n1176, C => 
                           Inst_CLB_switch_matrix_ConfigBits_84_port, ZN => 
                           n1010);
   U953 : AOI21D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_29_port, A2
                           => IJ_BEG_11_port, B => n888, ZN => n1299);
   U954 : INVD16 port map( I => n1299, ZN => E1BEG(2));
   U955 : BUFFD16 port map( I => n1332, Z => W2BEG(9));
   U956 : INVD16 port map( I => n810, ZN => N2BEG(5));
   U957 : INVD16 port map( I => n812, ZN => N2BEG(4));
   U958 : INVD16 port map( I => n814, ZN => N4BEG(7));
   U959 : INVD16 port map( I => n816, ZN => N4BEG(6));
   U960 : INVD16 port map( I => n818, ZN => E1BEG(1));
   U961 : INVD16 port map( I => n820, ZN => E1BEG(0));
   U962 : INVD16 port map( I => n822, ZN => E2BEG(7));
   U963 : INVD16 port map( I => n824, ZN => E2BEG(6));
   U964 : INVD16 port map( I => n826, ZN => E2BEG(5));
   U965 : INVD16 port map( I => n828, ZN => S1BEG(4));
   U966 : INVD16 port map( I => n830, ZN => S1BEG(3));
   U967 : INVD16 port map( I => n832, ZN => S1BEG(2));
   U968 : INVD16 port map( I => n834, ZN => S1BEG(1));
   U969 : INVD16 port map( I => n836, ZN => S1BEG(0));
   U970 : INVD16 port map( I => n838, ZN => S2BEG(7));
   U971 : INVD16 port map( I => n840, ZN => S2BEG(6));
   U972 : INVD16 port map( I => n842, ZN => S2BEG(5));
   U973 : INVD16 port map( I => n844, ZN => W1BEG(1));
   U974 : INVD16 port map( I => n846, ZN => W1BEG(0));
   U975 : INVD16 port map( I => n848, ZN => W2BEG(8));
   U976 : INVD16 port map( I => n850, ZN => W2BEG(7));
   U977 : INVD16 port map( I => n852, ZN => E2BEG(4));
   U978 : INVD16 port map( I => n854, ZN => S2BEG(9));
   U979 : INVD0 port map( I => n1342, ZN => n856);
   U980 : INVD0 port map( I => n856, ZN => n857);
   U981 : INVD16 port map( I => n856, ZN => CONFout);
   U982 : INVD0 port map( I => IJ_BEG_0_port, ZN => n464);
   U983 : INVD0 port map( I => IJ_BEG_10_port, ZN => n203);
   U984 : MAOI22D0 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_165_port, 
                           A2 => n526, B1 => OJ_BEG_2_port, B2 => 
                           Inst_CLB_switch_matrix_ConfigBits_165_port, ZN => 
                           n879);
   U985 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_158_port, 
                           A2 => n513, B1 => n906, B2 => n1102, ZN => 
                           IJ_BEG_4_port);
   U986 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_161_port, 
                           A2 => n138, B1 => n137, B2 => n136, ZN => n881);
   U987 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_15_port, ZN =>
                           n1243);
   U988 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_27_port, ZN =>
                           n1231);
   U989 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_82_port, ZN =>
                           n1176);
   U990 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_97_port, ZN =>
                           n1161);
   U991 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_115_port, ZN 
                           => n1143);
   U992 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_146_port, ZN 
                           => n1112);
   U993 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_153_port, ZN 
                           => n121);
   U994 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_171_port, ZN 
                           => n127);
   U995 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_C_values_10_port, ZN 
                           => n1065);
   U996 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_C_values_2_port, ZN =>
                           n1057);
   U997 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_102_port, ZN 
                           => n1156);
   U998 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_79_port, ZN =>
                           n1179);
   U999 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_62_port, ZN =>
                           n1196);
   U1000 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_74_port, ZN 
                           => n1184);
   U1001 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_54_port, ZN 
                           => n1204);
   U1002 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_38_port, ZN 
                           => n1220);
   U1003 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_16_port, ZN 
                           => n1242);
   U1004 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_10_port, ZN 
                           => n1248);
   U1005 : BUFFD16 port map( I => W2END(6), Z => W2BEG(0));
   U1006 : BUFFD16 port map( I => W2END(7), Z => W2BEG(1));
   U1007 : BUFFD16 port map( I => W2END(8), Z => W2BEG(2));
   U1008 : BUFFD16 port map( I => W2END(9), Z => W2BEG(3));
   U1009 : BUFFD16 port map( I => W2END(10), Z => W2BEG(4));
   U1010 : BUFFD16 port map( I => W2END(11), Z => W2BEG(5));
   U1011 : BUFFD16 port map( I => S2END(5), Z => S2BEG(0));
   U1012 : BUFFD16 port map( I => S2END(6), Z => S2BEG(1));
   U1013 : BUFFD16 port map( I => S2END(7), Z => S2BEG(2));
   U1014 : BUFFD16 port map( I => S2END(8), Z => S2BEG(3));
   U1015 : BUFFD16 port map( I => S2END(9), Z => S2BEG(4));
   U1016 : BUFFD16 port map( I => E2END(4), Z => E2BEG(0));
   U1017 : BUFFD16 port map( I => E2END(5), Z => E2BEG(1));
   U1018 : BUFFD16 port map( I => E2END(6), Z => E2BEG(2));
   U1019 : BUFFD16 port map( I => E2END(7), Z => E2BEG(3));
   U1020 : BUFFD16 port map( I => N4END(2), Z => N4BEG(0));
   U1021 : BUFFD16 port map( I => N4END(3), Z => N4BEG(1));
   U1022 : BUFFD16 port map( I => N4END(4), Z => N4BEG(2));
   U1023 : BUFFD16 port map( I => N4END(5), Z => N4BEG(3));
   U1024 : BUFFD16 port map( I => N4END(6), Z => N4BEG(4));
   U1025 : BUFFD16 port map( I => N4END(7), Z => N4BEG(5));
   U1026 : BUFFD16 port map( I => N2END(3), Z => N2BEG(0));
   U1027 : BUFFD16 port map( I => N2END(4), Z => N2BEG(1));
   U1028 : BUFFD16 port map( I => N2END(5), Z => N2BEG(2));
   U1029 : MUX4ND0 port map( I0 => Inst_clb_slice_4xLUT4_LUT_D_values_0_port, 
                           I1 => Inst_clb_slice_4xLUT4_LUT_D_values_1_port, I2 
                           => Inst_clb_slice_4xLUT4_LUT_D_values_2_port, I3 => 
                           Inst_clb_slice_4xLUT4_LUT_D_values_3_port, S0 => D0,
                           S1 => D1, ZN => n874);
   U1030 : INVD0 port map( I => D0, ZN => n868);
   U1031 : INVD0 port map( I => D1, ZN => n867);
   U1032 : AOI221D1 port map( A1 => D0, A2 => 
                           Inst_clb_slice_4xLUT4_LUT_D_values_11_port, B1 => 
                           n868, B2 => 
                           Inst_clb_slice_4xLUT4_LUT_D_values_10_port, C => 
                           n867, ZN => n864);
   U1033 : AOI221D1 port map( A1 => D0, A2 => 
                           Inst_clb_slice_4xLUT4_LUT_D_values_9_port, B1 => 
                           n868, B2 => 
                           Inst_clb_slice_4xLUT4_LUT_D_values_8_port, C => D1, 
                           ZN => n863);
   U1034 : AOI221D1 port map( A1 => D0, A2 => 
                           Inst_clb_slice_4xLUT4_LUT_D_values_7_port, B1 => 
                           n868, B2 => 
                           Inst_clb_slice_4xLUT4_LUT_D_values_6_port, C => n867
                           , ZN => n866);
   U1035 : AOI221D1 port map( A1 => D0, A2 => 
                           Inst_clb_slice_4xLUT4_LUT_D_values_5_port, B1 => 
                           n868, B2 => 
                           Inst_clb_slice_4xLUT4_LUT_D_values_4_port, C => D1, 
                           ZN => n865);
   U1036 : AOI221D1 port map( A1 => D0, A2 => conf_data_1_port, B1 => n868, B2 
                           => Inst_clb_slice_4xLUT4_LUT_D_values_14_port, C => 
                           n867, ZN => n870);
   U1037 : AOI221D1 port map( A1 => D0, A2 => 
                           Inst_clb_slice_4xLUT4_LUT_D_values_13_port, B1 => 
                           n868, B2 => 
                           Inst_clb_slice_4xLUT4_LUT_D_values_12_port, C => D1,
                           ZN => n869);
   U1038 : MUX4ND0 port map( I0 => n874, I1 => n873, I2 => n872, I3 => n871, S0
                           => D3, S1 => D2, ZN => D);
   U1039 : INVD0 port map( I => D, ZN => n506);
   U1040 : MUX4ND0 port map( I0 => n129, I1 => n130, I2 => n126, I3 => 
                           IJ_BEG_12_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_173_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_172_port, ZN => 
                           n526);
   U1041 : INVD0 port map( I => n526, ZN => IJ_BEG_9_port);
   U1042 : MUX4ND0 port map( I0 => IJ_BEG_9_port, I1 => IJ_BEG_10_port, I2 => 
                           IJ_BEG_11_port, I3 => IJ_BEG_12_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_149_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_150_port, ZN => 
                           n517);
   U1043 : MUX4ND0 port map( I0 => OJ_BEG_0_port, I1 => IJ_BEG_11_port, I2 => 
                           IJ_BEG_12_port, I3 => IJ_BEG_10_port, S0 => n1106, 
                           S1 => n1107, ZN => n518);
   U1044 : INVD0 port map( I => n517, ZN => n1011);
   U1045 : INVD0 port map( I => n518, ZN => n1015);
   U1046 : MUX4ND0 port map( I0 => TestOut, I1 => IJ_BEG_0_port, I2 => n1011, 
                           I3 => n1015, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_168_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_169_port, ZN => 
                           n876);
   U1047 : MUX4ND0 port map( I0 => IJ_BEG_9_port, I1 => IJ_BEG_11_port, I2 => 
                           IJ_BEG_10_port, I3 => IJ_BEG_12_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_169_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_168_port, ZN => 
                           n875);
   U1048 : MUX2ND0 port map( I0 => n876, I1 => n875, S => 
                           Inst_CLB_switch_matrix_ConfigBits_170_port, ZN => 
                           IJ_BEG_8_port);
   U1049 : INVD0 port map( I => IJ_BEG_8_port, ZN => n529);
   U1050 : INVD0 port map( I => TestOut, ZN => n893);
   U1051 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_165_port, 
                           A2 => n893, B1 => n507, B2 => n1097, ZN => n880);
   U1052 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_165_port, 
                           A2 => n517, B1 => n464, B2 => n1097, ZN => n878);
   U1053 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_165_port, 
                           A2 => n218, B1 => n203, B2 => n1097, ZN => n877);
   U1054 : MUX4ND0 port map( I0 => n880, I1 => n879, I2 => n878, I3 => n877, S0
                           => Inst_CLB_switch_matrix_ConfigBits_167_port, S1 =>
                           Inst_CLB_switch_matrix_ConfigBits_166_port, ZN => 
                           n270);
   U1055 : INVD0 port map( I => n270, ZN => IJ_BEG_7_port);
   U1056 : MUX2ND0 port map( I0 => n881, I1 => n140, S => 
                           Inst_CLB_switch_matrix_ConfigBits_160_port, ZN => 
                           n528);
   U1057 : INVD0 port map( I => n528, ZN => IJ_BEG_5_port);
   U1058 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_180_port, 
                           A2 => n203, B1 => n270, B2 => n1088, ZN => 
                           OJ_BEG_1_port);
   U1059 : MUX4ND0 port map( I0 => D, I1 => DQ, I2 => TestOut, I3 => 
                           IJ_BEG_0_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_162_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_163_port, ZN => 
                           n883);
   U1060 : MUX2ND0 port map( I0 => n883, I1 => n882, S => 
                           Inst_CLB_switch_matrix_ConfigBits_164_port, ZN => 
                           IJ_BEG_6_port);
   U1061 : MUX4ND0 port map( I0 => E1END(1), I1 => IJ_BEG_7_port, I2 => 
                           E1END(2), I3 => IJ_BEG_8_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_19_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_17_port, ZN => 
                           n885);
   U1062 : MUX4ND0 port map( I0 => N4END(1), I1 => IJ_BEG_5_port, I2 => 
                           E1END(0), I3 => IJ_BEG_6_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_19_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_17_port, ZN => 
                           n884);
   U1063 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_18_port, ZN 
                           => n1240);
   U1064 : MUX4ND0 port map( I0 => E2END(0), I1 => IJ_BEG_9_port, I2 => 
                           E2END(1), I3 => IJ_BEG_10_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_28_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_26_port, ZN => 
                           n887);
   U1065 : MUX4ND0 port map( I0 => E1END(2), I1 => DQ, I2 => E1END(3), I3 => 
                           IJ_BEG_8_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_28_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_26_port, ZN => 
                           n886);
   U1066 : MUX4ND0 port map( I0 => E1END(2), I1 => IJ_BEG_8_port, I2 => 
                           E1END(3), I3 => IJ_BEG_9_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_22_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_20_port, ZN => 
                           n890);
   U1067 : MUX4ND0 port map( I0 => E1END(0), I1 => IJ_BEG_6_port, I2 => 
                           E1END(1), I3 => IJ_BEG_7_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_22_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_20_port, ZN => 
                           n889);
   U1068 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_21_port, ZN 
                           => n1237);
   U1069 : MUX4ND0 port map( I0 => E2END(3), I1 => IJ_BEG_0_port, I2 => 
                           S1END(0), I3 => n1011, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_39_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_37_port, ZN => 
                           n892);
   U1070 : MUX4ND0 port map( I0 => E2END(1), I1 => DQ, I2 => E2END(2), I3 => 
                           TestOut, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_39_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_37_port, ZN => 
                           n891);
   U1071 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_34_port, ZN 
                           => n1224);
   U1072 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_34_port, 
                           A2 => n893, B1 => n507, B2 => n1224, ZN => n894);
   U1073 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_35_port, ZN 
                           => n1223);
   U1074 : MUX4ND0 port map( I0 => E2END(0), I1 => E2END(2), I2 => E2END(1), I3
                           => E2END(3), S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_35_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_34_port, ZN => 
                           n895);
   U1075 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_36_port, ZN 
                           => n1222);
   U1076 : MUX4ND0 port map( I0 => W1END(5), I1 => TestOut, I2 => W2END(0), I3 
                           => IJ_BEG_0_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_95_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_93_port, ZN => 
                           n900);
   U1077 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_93_port, ZN 
                           => n1165);
   U1078 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_93_port, 
                           A2 => IJ_BEG_11_port, B1 => IJ_BEG_10_port, B2 => 
                           n1165, ZN => n899);
   U1079 : MUX4ND0 port map( I0 => W2END(1), I1 => n1011, I2 => W2END(2), I3 =>
                           n1015, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_95_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_93_port, ZN => 
                           n898);
   U1080 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_93_port, 
                           A2 => OJ_BEG_0_port, B1 => IJ_BEG_12_port, B2 => 
                           n1165, ZN => n897);
   U1081 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_153_port, 
                           A2 => OJ_BEG_0_port, B1 => IJ_BEG_12_port, B2 => 
                           n121, ZN => n901);
   U1082 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_154_port, 
                           A2 => n901, B1 => n123, B2 => n1105, ZN => n902);
   U1083 : MUX2ND0 port map( I0 => n902, I1 => OJ_BEG_1_port, S => 
                           Inst_CLB_switch_matrix_ConfigBits_155_port, ZN => 
                           n514);
   U1084 : INVD0 port map( I => n514, ZN => IJ_BEG_3_port);
   U1085 : MUX4ND0 port map( I0 => S2END(0), I1 => n1015, I2 => S2END(1), I3 =>
                           IJ_BEG_3_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_57_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_55_port, ZN => 
                           n904);
   U1086 : MUX4ND0 port map( I0 => S1END(3), I1 => IJ_BEG_0_port, I2 => 
                           S1END(4), I3 => n1011, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_57_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_55_port, ZN => 
                           n903);
   U1087 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_56_port, ZN 
                           => n1202);
   U1088 : INVD0 port map( I => IJ_BEG_12_port, ZN => n993);
   U1089 : MAOI22D0 port map( A1 => n993, A2 => n505, B1 => n505, B2 => 
                           OJ_BEG_0_port, ZN => n905);
   U1090 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_157_port, 
                           A2 => n905, B1 => n509, B2 => n1103, ZN => n906);
   U1091 : MUX4ND0 port map( I0 => n1011, I1 => n1015, I2 => IJ_BEG_3_port, I3 
                           => IJ_BEG_4_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_133_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_134_port, ZN => 
                           n907);
   U1092 : MUX4ND0 port map( I0 => TestOut, I1 => IJ_BEG_0_port, I2 => n1011, 
                           I3 => n1015, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_129_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_130_port, ZN => 
                           n908);
   U1093 : NR2D0 port map( A1 => n907, A2 => n908, ZN => n926);
   U1094 : CKND2D0 port map( A1 => n907, A2 => n908, ZN => n918);
   U1095 : INVD0 port map( I => n907, ZN => n909);
   U1096 : CKND2D0 port map( A1 => n909, A2 => n908, ZN => n923);
   U1097 : INVD0 port map( I => n923, ZN => n915);
   U1098 : MUX4ND0 port map( I0 => IJ_BEG_0_port, I1 => n1015, I2 => n1011, I3 
                           => IJ_BEG_3_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_132_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_131_port, ZN => 
                           n922);
   U1099 : AOI21D1 port map( A1 => Inst_clb_slice_4xLUT4_LUT_C_values_14_port, 
                           A2 => n915, B => n922, ZN => n911);
   U1100 : NR2D0 port map( A1 => n909, A2 => n908, ZN => n919);
   U1101 : AOI22D1 port map( A1 => Inst_clb_slice_4xLUT4_LUT_C_values_15_port, 
                           A2 => n926, B1 => 
                           Inst_clb_slice_4xLUT4_LUT_C_values_11_port, B2 => 
                           n919, ZN => n910);
   U1102 : OAI211D1 port map( A1 => n1065, A2 => n918, B => n911, C => n910, ZN
                           => n914);
   U1103 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_C_values_12_port, ZN 
                           => n1067);
   U1104 : INVD0 port map( I => n918, ZN => n920);
   U1105 : AOI22D1 port map( A1 => n920, A2 => 
                           Inst_clb_slice_4xLUT4_LUT_C_values_8_port, B1 => 
                           n919, B2 => 
                           Inst_clb_slice_4xLUT4_LUT_C_values_9_port, ZN => 
                           n912);
   U1106 : OAI211D1 port map( A1 => n1067, A2 => n923, B => n922, C => n912, ZN
                           => n913);
   U1107 : AOI32D1 port map( A1 => n926, A2 => n914, A3 => 
                           Inst_clb_slice_4xLUT4_LUT_C_values_13_port, B1 => 
                           n913, B2 => n914, ZN => n929);
   U1108 : AOI21D1 port map( A1 => n915, A2 => 
                           Inst_clb_slice_4xLUT4_LUT_C_values_6_port, B => n922
                           , ZN => n917);
   U1109 : AOI22D1 port map( A1 => n926, A2 => 
                           Inst_clb_slice_4xLUT4_LUT_C_values_7_port, B1 => 
                           n919, B2 => 
                           Inst_clb_slice_4xLUT4_LUT_C_values_3_port, ZN => 
                           n916);
   U1110 : OAI211D1 port map( A1 => n918, A2 => n1057, B => n917, C => n916, ZN
                           => n925);
   U1111 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_C_values_4_port, ZN 
                           => n1059);
   U1112 : AOI22D1 port map( A1 => n920, A2 => 
                           Inst_clb_slice_4xLUT4_LUT_C_values_0_port, B1 => 
                           n919, B2 => 
                           Inst_clb_slice_4xLUT4_LUT_C_values_1_port, ZN => 
                           n921);
   U1113 : OAI211D1 port map( A1 => n1059, A2 => n923, B => n922, C => n921, ZN
                           => n924);
   U1114 : AOI32D1 port map( A1 => n926, A2 => n925, A3 => 
                           Inst_clb_slice_4xLUT4_LUT_C_values_5_port, B1 => 
                           n924, B2 => n925, ZN => n928);
   U1115 : MUX4ND0 port map( I0 => n1015, I1 => IJ_BEG_4_port, I2 => 
                           IJ_BEG_3_port, I3 => IJ_BEG_5_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_136_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_135_port, ZN => 
                           n927);
   U1116 : MUX2ND0 port map( I0 => n929, I1 => n928, S => n927, ZN => C);
   U1117 : MUX4ND0 port map( I0 => D, I1 => TestOut, I2 => DQ, I3 => 
                           IJ_BEG_0_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_126_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_125_port, ZN => 
                           n930);
   U1118 : MUX4ND0 port map( I0 => C, I1 => CQ, I2 => D, I3 => DQ, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_121_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_122_port, ZN => 
                           n931);
   U1119 : NR2D0 port map( A1 => n930, A2 => n931, ZN => n948);
   U1120 : CKND2D0 port map( A1 => n930, A2 => n931, ZN => n941);
   U1121 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_B_values_10_port, ZN 
                           => n1049);
   U1122 : INVD0 port map( I => n930, ZN => n932);
   U1123 : CKND2D0 port map( A1 => n932, A2 => n931, ZN => n946);
   U1124 : INVD0 port map( I => n946, ZN => n938);
   U1125 : MUX4ND0 port map( I0 => CQ, I1 => D, I2 => DQ, I3 => TestOut, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_123_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_124_port, ZN => 
                           n944);
   U1126 : AOI21D1 port map( A1 => n938, A2 => 
                           Inst_clb_slice_4xLUT4_LUT_B_values_14_port, B => 
                           n944, ZN => n934);
   U1127 : NR2D0 port map( A1 => n932, A2 => n931, ZN => n942);
   U1128 : AOI22D1 port map( A1 => n948, A2 => 
                           Inst_clb_slice_4xLUT4_LUT_B_values_15_port, B1 => 
                           n942, B2 => 
                           Inst_clb_slice_4xLUT4_LUT_B_values_11_port, ZN => 
                           n933);
   U1129 : OAI211D1 port map( A1 => n941, A2 => n1049, B => n934, C => n933, ZN
                           => n937);
   U1130 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_B_values_12_port, ZN 
                           => n1051);
   U1131 : INVD0 port map( I => n941, ZN => n943);
   U1132 : AOI22D1 port map( A1 => Inst_clb_slice_4xLUT4_LUT_B_values_8_port, 
                           A2 => n943, B1 => 
                           Inst_clb_slice_4xLUT4_LUT_B_values_9_port, B2 => 
                           n942, ZN => n935);
   U1133 : OAI211D1 port map( A1 => n1051, A2 => n946, B => n935, C => n944, ZN
                           => n936);
   U1134 : AOI32D1 port map( A1 => n948, A2 => n937, A3 => 
                           Inst_clb_slice_4xLUT4_LUT_B_values_13_port, B1 => 
                           n936, B2 => n937, ZN => n952);
   U1135 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_B_values_2_port, ZN 
                           => n1041);
   U1136 : AOI21D1 port map( A1 => n938, A2 => 
                           Inst_clb_slice_4xLUT4_LUT_B_values_6_port, B => n944
                           , ZN => n940);
   U1137 : AOI22D1 port map( A1 => n948, A2 => 
                           Inst_clb_slice_4xLUT4_LUT_B_values_7_port, B1 => 
                           n942, B2 => 
                           Inst_clb_slice_4xLUT4_LUT_B_values_3_port, ZN => 
                           n939);
   U1138 : OAI211D1 port map( A1 => n941, A2 => n1041, B => n940, C => n939, ZN
                           => n949);
   U1139 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_B_values_4_port, ZN 
                           => n1043);
   U1140 : AOI22D1 port map( A1 => n943, A2 => 
                           Inst_clb_slice_4xLUT4_LUT_B_values_0_port, B1 => 
                           n942, B2 => 
                           Inst_clb_slice_4xLUT4_LUT_B_values_1_port, ZN => 
                           n945);
   U1141 : OAI211D1 port map( A1 => n946, A2 => n1043, B => n945, C => n944, ZN
                           => n947);
   U1142 : AOI32D1 port map( A1 => Inst_clb_slice_4xLUT4_LUT_B_values_5_port, 
                           A2 => n949, A3 => n948, B1 => n947, B2 => n949, ZN 
                           => n951);
   U1143 : MUX4ND0 port map( I0 => DQ, I1 => IJ_BEG_0_port, I2 => TestOut, I3 
                           => n1011, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_128_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_127_port, ZN => 
                           n950);
   U1144 : MUX2ND0 port map( I0 => n952, I1 => n951, S => n950, ZN => B);
   U1145 : MUX4ND0 port map( I0 => C, I1 => BQ, I2 => B, I3 => AQ, S0 => n1143,
                           S1 => n1142, ZN => n958);
   U1146 : INVD0 port map( I => n958, ZN => n959);
   U1147 : MUX4ND0 port map( I0 => Inst_clb_slice_4xLUT4_LUT_A_values_0_port, 
                           I1 => Inst_clb_slice_4xLUT4_LUT_A_values_1_port, I2 
                           => Inst_clb_slice_4xLUT4_LUT_A_values_2_port, I3 => 
                           Inst_clb_slice_4xLUT4_LUT_A_values_3_port, S0 => A0,
                           S1 => n959, ZN => n967);
   U1148 : INVD0 port map( I => A0, ZN => n957);
   U1149 : AOI221D1 port map( A1 => n959, A2 => 
                           Inst_clb_slice_4xLUT4_LUT_A_values_11_port, B1 => 
                           n958, B2 => 
                           Inst_clb_slice_4xLUT4_LUT_A_values_9_port, C => n957
                           , ZN => n954);
   U1150 : AOI221D1 port map( A1 => n959, A2 => 
                           Inst_clb_slice_4xLUT4_LUT_A_values_10_port, B1 => 
                           n958, B2 => 
                           Inst_clb_slice_4xLUT4_LUT_A_values_8_port, C => A0, 
                           ZN => n953);
   U1151 : AOI221D1 port map( A1 => n959, A2 => 
                           Inst_clb_slice_4xLUT4_LUT_A_values_7_port, B1 => 
                           n958, B2 => 
                           Inst_clb_slice_4xLUT4_LUT_A_values_5_port, C => n957
                           , ZN => n956);
   U1152 : AOI221D1 port map( A1 => n959, A2 => 
                           Inst_clb_slice_4xLUT4_LUT_A_values_6_port, B1 => 
                           n958, B2 => 
                           Inst_clb_slice_4xLUT4_LUT_A_values_4_port, C => A0, 
                           ZN => n955);
   U1153 : AOI221D1 port map( A1 => n959, A2 => 
                           Inst_clb_slice_4xLUT4_LUT_A_values_15_port, B1 => 
                           n958, B2 => 
                           Inst_clb_slice_4xLUT4_LUT_A_values_13_port, C => 
                           n957, ZN => n961);
   U1154 : AOI221D1 port map( A1 => n959, A2 => 
                           Inst_clb_slice_4xLUT4_LUT_A_values_14_port, B1 => 
                           n958, B2 => 
                           Inst_clb_slice_4xLUT4_LUT_A_values_12_port, C => A0,
                           ZN => n960);
   U1155 : OR2D1 port map( A1 => n961, A2 => n960, Z => n964);
   U1156 : MUX4D1 port map( I0 => BQ, I1 => C, I2 => CQ, I3 => D, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_119_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_120_port, Z => 
                           n963);
   U1157 : MUX4D1 port map( I0 => B, I1 => C, I2 => BQ, I3 => CQ, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_118_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_117_port, Z => 
                           n962);
   U1158 : MUX4ND0 port map( I0 => n967, I1 => n966, I2 => n965, I3 => n964, S0
                           => n963, S1 => n962, ZN => A);
   U1159 : MUX4D1 port map( I0 => W2END(5), I1 => AQ, I2 => A, I3 => B, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_112_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_111_port, Z => 
                           n1330);
   U1160 : MUX4ND0 port map( I0 => S1END(3), I1 => IJ_BEG_4_port, I2 => 
                           S1END(4), I3 => IJ_BEG_5_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_51_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_49_port, ZN => 
                           n969);
   U1161 : MUX4ND0 port map( I0 => S1END(1), I1 => n1015, I2 => S1END(2), I3 =>
                           IJ_BEG_3_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_51_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_49_port, ZN => 
                           n968);
   U1162 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_50_port, ZN 
                           => n1208);
   U1163 : MUX4ND0 port map( I0 => S1END(1), I1 => n1015, I2 => S1END(2), I3 =>
                           IJ_BEG_3_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_45_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_43_port, ZN => 
                           n971);
   U1164 : MUX4ND0 port map( I0 => E2END(3), I1 => IJ_BEG_0_port, I2 => 
                           S1END(0), I3 => n1011, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_45_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_43_port, ZN => 
                           n970);
   U1165 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_44_port, ZN 
                           => n1214);
   U1166 : MUX4ND0 port map( I0 => S1END(2), I1 => IJ_BEG_3_port, I2 => 
                           S1END(3), I3 => IJ_BEG_4_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_48_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_46_port, ZN => 
                           n973);
   U1167 : MUX4ND0 port map( I0 => S1END(0), I1 => n1011, I2 => S1END(1), I3 =>
                           n1015, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_48_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_46_port, ZN => 
                           n972);
   U1168 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_47_port, ZN 
                           => n1211);
   U1169 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_11_port, ZN 
                           => n1247);
   U1170 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_11_port, 
                           A2 => IJ_BEG_6_port, B1 => IJ_BEG_5_port, B2 => 
                           n1247, ZN => n975);
   U1171 : MUX4ND0 port map( I0 => N2END(2), I1 => N4END(1), I2 => N4END(0), I3
                           => E1END(0), S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_12_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_11_port, ZN => 
                           n974);
   U1172 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_13_port, ZN 
                           => n1245);
   U1173 : MUX4ND0 port map( I0 => W2END(4), I1 => IJ_BEG_4_port, I2 => 
                           W2END(5), I3 => IJ_BEG_5_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_106_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_104_port, ZN => 
                           n977);
   U1174 : MUX4ND0 port map( I0 => W2END(2), I1 => n1015, I2 => W2END(3), I3 =>
                           IJ_BEG_3_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_106_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_104_port, ZN => 
                           n976);
   U1175 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_105_port, ZN 
                           => n1153);
   U1176 : MUX4ND0 port map( I0 => S2END(3), I1 => IJ_BEG_5_port, I2 => 
                           S2END(4), I3 => IJ_BEG_6_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_66_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_64_port, ZN => 
                           n979);
   U1177 : MUX4ND0 port map( I0 => S2END(1), I1 => IJ_BEG_3_port, I2 => 
                           S2END(2), I3 => IJ_BEG_4_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_66_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_64_port, ZN => 
                           n978);
   U1178 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_65_port, ZN 
                           => n1193);
   U1179 : MUX4ND0 port map( I0 => W2END(3), I1 => IJ_BEG_3_port, I2 => 
                           W2END(4), I3 => IJ_BEG_4_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_103_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_101_port, ZN => 
                           n981);
   U1180 : MUX4ND0 port map( I0 => W2END(1), I1 => n1011, I2 => W2END(2), I3 =>
                           n1015, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_103_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_101_port, ZN => 
                           n980);
   U1181 : MUX4ND0 port map( I0 => W2END(0), I1 => IJ_BEG_0_port, I2 => 
                           W2END(1), I3 => n1011, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_99_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_97_port, ZN => 
                           n985);
   U1182 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_97_port, 
                           A2 => IJ_BEG_12_port, B1 => IJ_BEG_11_port, B2 => 
                           n1161, ZN => n984);
   U1183 : MUX4ND0 port map( I0 => W2END(2), I1 => n1015, I2 => W2END(3), I3 =>
                           IJ_BEG_3_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_99_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_97_port, ZN => 
                           n983);
   U1184 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_97_port, 
                           A2 => OJ_BEG_1_port, B1 => OJ_BEG_0_port, B2 => 
                           n1161, ZN => n982);
   U1185 : MUX4ND0 port map( I0 => N2END(1), I1 => N4END(0), I2 => N2END(2), I3
                           => N4END(1), S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_9_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_8_port, ZN => n986
                           );
   U1186 : MUX4ND0 port map( I0 => S2END(4), I1 => IJ_BEG_6_port, I2 => 
                           W1END(0), I3 => IJ_BEG_7_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_69_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_67_port, ZN => 
                           n988);
   U1187 : MUX4ND0 port map( I0 => S2END(2), I1 => IJ_BEG_4_port, I2 => 
                           S2END(3), I3 => IJ_BEG_5_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_69_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_67_port, ZN => 
                           n987);
   U1188 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_68_port, ZN 
                           => n1190);
   U1189 : MUX4ND0 port map( I0 => W1END(4), I1 => DQ, I2 => W1END(5), I3 => 
                           TestOut, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_91_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_89_port, ZN => 
                           n992);
   U1190 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_89_port, ZN 
                           => n1169);
   U1191 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_89_port, 
                           A2 => IJ_BEG_10_port, B1 => IJ_BEG_9_port, B2 => 
                           n1169, ZN => n991);
   U1192 : MUX4ND0 port map( I0 => W2END(0), I1 => IJ_BEG_0_port, I2 => 
                           W2END(1), I3 => n1011, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_91_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_89_port, ZN => 
                           n990);
   U1193 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_89_port, 
                           A2 => IJ_BEG_12_port, B1 => IJ_BEG_11_port, B2 => 
                           n1169, ZN => n989);
   U1194 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_30_port, ZN 
                           => n1228);
   U1195 : MUX4ND0 port map( I0 => E2END(1), I1 => IJ_BEG_9_port, I2 => 
                           E2END(2), I3 => IJ_BEG_10_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_32_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_30_port, ZN => 
                           n995);
   U1196 : MUX4ND0 port map( I0 => E1END(3), I1 => DQ, I2 => E2END(0), I3 => 
                           TestOut, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_32_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_30_port, ZN => 
                           n994);
   U1197 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_31_port, ZN 
                           => n1227);
   U1198 : MUX4ND0 port map( I0 => S2END(2), I1 => IJ_BEG_4_port, I2 => 
                           S2END(3), I3 => IJ_BEG_5_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_63_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_61_port, ZN => 
                           n998);
   U1199 : MUX4ND0 port map( I0 => S2END(0), I1 => n1015, I2 => S2END(1), I3 =>
                           IJ_BEG_3_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_63_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_61_port, ZN => 
                           n997);
   U1200 : MUX4ND0 port map( I0 => E1END(3), I1 => IJ_BEG_9_port, I2 => 
                           E2END(0), I3 => IJ_BEG_10_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_25_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_23_port, ZN => 
                           n1000);
   U1201 : MUX4ND0 port map( I0 => E1END(1), I1 => IJ_BEG_7_port, I2 => 
                           E1END(2), I3 => IJ_BEG_8_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_25_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_23_port, ZN => 
                           n999);
   U1202 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_24_port, ZN 
                           => n1234);
   U1203 : MUX4ND0 port map( I0 => S2END(4), I1 => W1END(1), I2 => W1END(0), I3
                           => W1END(2), S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_73_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_72_port, ZN => 
                           n1001);
   U1204 : MUX4ND0 port map( I0 => W1END(3), I1 => IJ_BEG_8_port, I2 => 
                           W1END(4), I3 => IJ_BEG_9_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_80_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_78_port, ZN => 
                           n1003);
   U1205 : MUX4ND0 port map( I0 => W1END(1), I1 => DQ, I2 => W1END(2), I3 => 
                           IJ_BEG_7_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_80_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_78_port, ZN => 
                           n1002);
   U1206 : MUX4ND0 port map( I0 => S1END(0), I1 => n1011, I2 => S1END(1), I3 =>
                           n1015, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_42_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_40_port, ZN => 
                           n1005);
   U1207 : MUX4ND0 port map( I0 => E2END(2), I1 => TestOut, I2 => E2END(3), I3 
                           => IJ_BEG_0_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_42_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_40_port, ZN => 
                           n1004);
   U1208 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_41_port, ZN 
                           => n1217);
   U1209 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_75_port, ZN 
                           => n1183);
   U1210 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_75_port, 
                           A2 => IJ_BEG_8_port, B1 => IJ_BEG_7_port, B2 => 
                           n1183, ZN => n1007);
   U1211 : MUX4ND0 port map( I0 => W1END(0), I1 => W1END(2), I2 => W1END(1), I3
                           => W1END(3), S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_76_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_75_port, ZN => 
                           n1006);
   U1212 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_77_port, ZN 
                           => n1181);
   U1213 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_81_port, ZN 
                           => n1177);
   U1214 : MUX4ND0 port map( I0 => W1END(4), I1 => IJ_BEG_7_port, I2 => 
                           W1END(5), I3 => IJ_BEG_8_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_83_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_81_port, ZN => 
                           n1009);
   U1215 : MUX4ND0 port map( I0 => W1END(2), I1 => DQ, I2 => W1END(3), I3 => 
                           TestOut, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_83_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_81_port, ZN => 
                           n1008);
   U1216 : MUX4ND0 port map( I0 => S2END(1), I1 => IJ_BEG_3_port, I2 => 
                           S2END(2), I3 => IJ_BEG_4_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_60_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_58_port, ZN => 
                           n1013);
   U1217 : MUX4ND0 port map( I0 => S1END(4), I1 => n1011, I2 => S2END(0), I3 =>
                           n1015, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_60_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_58_port, ZN => 
                           n1012);
   U1218 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_59_port, ZN 
                           => n1199);
   U1219 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_52_port, ZN 
                           => n1206);
   U1220 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_52_port, 
                           A2 => n517, B1 => n464, B2 => n1206, ZN => n1014);
   U1221 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_53_port, ZN 
                           => n1205);
   U1222 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_53_port, 
                           A2 => n1015, B1 => n1014, B2 => n1205, ZN => n1017);
   U1223 : MUX4ND0 port map( I0 => S1END(2), I1 => S1END(4), I2 => S1END(3), I3
                           => S2END(0), S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_53_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_52_port, ZN => 
                           n1016);
   U1224 : MUX4D1 port map( I0 => W2END(4), I1 => A, I2 => W2END(5), I3 => AQ, 
                           S0 => Inst_CLB_switch_matrix_ConfigBits_110_port, S1
                           => Inst_CLB_switch_matrix_ConfigBits_109_port, Z => 
                           n1331);
   U1225 : INVD0 port map( I => IJ_BEG_6_port, ZN => n525);
   U1226 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_14_port, ZN 
                           => n1244);
   U1227 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_14_port, 
                           A2 => n525, B1 => n528, B2 => n1244, ZN => n1018);
   U1228 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_15_port, 
                           A2 => IJ_BEG_7_port, B1 => n1018, B2 => n1243, ZN =>
                           n1020);
   U1229 : MUX4ND0 port map( I0 => N4END(0), I1 => E1END(0), I2 => N4END(1), I3
                           => E1END(1), S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_15_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_14_port, ZN => 
                           n1019);
   U1230 : MUX4ND0 port map( I0 => W1END(3), I1 => DQ, I2 => W1END(4), I3 => 
                           TestOut, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_87_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_85_port, ZN => 
                           n1023);
   U1231 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_85_port, ZN 
                           => n1173);
   U1232 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_85_port, 
                           A2 => IJ_BEG_10_port, B1 => IJ_BEG_9_port, B2 => 
                           n1173, ZN => n1022);
   U1233 : MUX4ND0 port map( I0 => W1END(5), I1 => IJ_BEG_0_port, I2 => 
                           W2END(0), I3 => IJ_BEG_8_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_87_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_85_port, ZN => 
                           n1021);
   U1234 : INVD0 port map( I => IJ_BEG_4_port, ZN => n515);
   U1235 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_A_values_1_port, ZN 
                           => n1024);
   U1236 : MAOI22D0 port map( A1 => n1024, A2 => n780, B1 => n781, B2 => 
                           Inst_clb_slice_4xLUT4_LUT_A_values_0_port, ZN => 
                           n775);
   U1237 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_1_port, ZN =>
                           n1256);
   U1238 : MAOI22D0 port map( A1 => MODE, A2 => n1256, B1 => 
                           Inst_CLB_switch_matrix_ConfigBits_0_port, B2 => MODE
                           , ZN => n530);
   U1239 : INVD0 port map( I => conf_data_2_port, ZN => n1086);
   U1240 : AOI22D1 port map( A1 => MODE, A2 => n1086, B1 => n856, B2 => n777, 
                           ZN => n711);
   U1241 : AOI22D1 port map( A1 => MODE, A2 => n856, B1 => n1088, B2 => n778, 
                           ZN => n710);
   U1242 : MUX4ND0 port map( I0 => n526, I1 => n270, I2 => n203, I3 => n529, S0
                           => n1112, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_145_port, ZN => 
                           TestIn);
   U1243 : AOI22D1 port map( A1 => Inst_CLB_switch_matrix_ConfigBits_175_port, 
                           A2 => n521, B1 => n520, B2 => n1089, ZN => n523);
   U1244 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_A_values_2_port, ZN 
                           => n1025);
   U1245 : AOI22D1 port map( A1 => MODE, A2 => n1024, B1 => n1025, B2 => n780, 
                           ZN => n774);
   U1246 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_A_values_3_port, ZN 
                           => n1026);
   U1247 : AOI22D1 port map( A1 => MODE, A2 => n1025, B1 => n1026, B2 => n782, 
                           ZN => n773);
   U1248 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_A_values_4_port, ZN 
                           => n1027);
   U1249 : AOI22D1 port map( A1 => MODE, A2 => n1026, B1 => n1027, B2 => n780, 
                           ZN => n772);
   U1250 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_A_values_5_port, ZN 
                           => n1028);
   U1251 : AOI22D1 port map( A1 => MODE, A2 => n1027, B1 => n1028, B2 => n780, 
                           ZN => n771);
   U1252 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_A_values_6_port, ZN 
                           => n1029);
   U1253 : AOI22D1 port map( A1 => MODE, A2 => n1028, B1 => n1029, B2 => n779, 
                           ZN => n770);
   U1254 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_A_values_7_port, ZN 
                           => n1030);
   U1255 : AOI22D1 port map( A1 => MODE, A2 => n1029, B1 => n1030, B2 => n777, 
                           ZN => n769);
   U1256 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_A_values_8_port, ZN 
                           => n1031);
   U1257 : AOI22D1 port map( A1 => MODE, A2 => n1030, B1 => n1031, B2 => n777, 
                           ZN => n768);
   U1258 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_A_values_9_port, ZN 
                           => n1032);
   U1259 : AOI22D1 port map( A1 => MODE, A2 => n1031, B1 => n1032, B2 => n777, 
                           ZN => n767);
   U1260 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_A_values_10_port, ZN 
                           => n1033);
   U1261 : AOI22D1 port map( A1 => MODE, A2 => n1032, B1 => n1033, B2 => n777, 
                           ZN => n766);
   U1262 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_A_values_11_port, ZN 
                           => n1034);
   U1263 : AOI22D1 port map( A1 => MODE, A2 => n1033, B1 => n1034, B2 => n777, 
                           ZN => n765);
   U1264 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_A_values_12_port, ZN 
                           => n1035);
   U1265 : AOI22D1 port map( A1 => MODE, A2 => n1034, B1 => n1035, B2 => n778, 
                           ZN => n764);
   U1266 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_A_values_13_port, ZN 
                           => n1036);
   U1267 : AOI22D1 port map( A1 => MODE, A2 => n1035, B1 => n1036, B2 => n782, 
                           ZN => n763);
   U1268 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_A_values_14_port, ZN 
                           => n1037);
   U1269 : AOI22D1 port map( A1 => MODE, A2 => n1036, B1 => n1037, B2 => n779, 
                           ZN => n762);
   U1270 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_A_values_15_port, ZN 
                           => n1038);
   U1271 : AOI22D1 port map( A1 => MODE, A2 => n1037, B1 => n1038, B2 => n777, 
                           ZN => n761);
   U1272 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_B_values_0_port, ZN 
                           => n1039);
   U1273 : AOI22D1 port map( A1 => MODE, A2 => n1038, B1 => n1039, B2 => n778, 
                           ZN => n760);
   U1274 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_B_values_1_port, ZN 
                           => n1040);
   U1275 : AOI22D1 port map( A1 => MODE, A2 => n1039, B1 => n1040, B2 => n778, 
                           ZN => n759);
   U1276 : AOI22D1 port map( A1 => MODE, A2 => n1040, B1 => n1041, B2 => n782, 
                           ZN => n758);
   U1277 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_B_values_3_port, ZN 
                           => n1042);
   U1278 : AOI22D1 port map( A1 => MODE, A2 => n1041, B1 => n1042, B2 => n778, 
                           ZN => n757);
   U1279 : AOI22D1 port map( A1 => MODE, A2 => n1042, B1 => n1043, B2 => n780, 
                           ZN => n756);
   U1280 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_B_values_5_port, ZN 
                           => n1044);
   U1281 : AOI22D1 port map( A1 => MODE, A2 => n1043, B1 => n1044, B2 => n778, 
                           ZN => n755);
   U1282 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_B_values_6_port, ZN 
                           => n1045);
   U1283 : AOI22D1 port map( A1 => MODE, A2 => n1044, B1 => n1045, B2 => n781, 
                           ZN => n754);
   U1284 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_B_values_7_port, ZN 
                           => n1046);
   U1285 : AOI22D1 port map( A1 => MODE, A2 => n1045, B1 => n1046, B2 => n781, 
                           ZN => n753);
   U1286 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_B_values_8_port, ZN 
                           => n1047);
   U1287 : AOI22D1 port map( A1 => MODE, A2 => n1046, B1 => n1047, B2 => n778, 
                           ZN => n752);
   U1288 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_B_values_9_port, ZN 
                           => n1048);
   U1289 : AOI22D1 port map( A1 => MODE, A2 => n1047, B1 => n1048, B2 => n778, 
                           ZN => n751);
   U1290 : AOI22D1 port map( A1 => MODE, A2 => n1048, B1 => n1049, B2 => n777, 
                           ZN => n750);
   U1291 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_B_values_11_port, ZN 
                           => n1050);
   U1292 : AOI22D1 port map( A1 => MODE, A2 => n1049, B1 => n1050, B2 => n777, 
                           ZN => n749);
   U1293 : AOI22D1 port map( A1 => MODE, A2 => n1050, B1 => n1051, B2 => n778, 
                           ZN => n748);
   U1294 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_B_values_13_port, ZN 
                           => n1052);
   U1295 : AOI22D1 port map( A1 => MODE, A2 => n1051, B1 => n1052, B2 => n778, 
                           ZN => n747);
   U1296 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_B_values_14_port, ZN 
                           => n1053);
   U1297 : AOI22D1 port map( A1 => MODE, A2 => n1052, B1 => n1053, B2 => n777, 
                           ZN => n746);
   U1298 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_B_values_15_port, ZN 
                           => n1054);
   U1299 : AOI22D1 port map( A1 => MODE, A2 => n1053, B1 => n1054, B2 => n777, 
                           ZN => n745);
   U1300 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_C_values_0_port, ZN 
                           => n1055);
   U1301 : AOI22D1 port map( A1 => MODE, A2 => n1054, B1 => n1055, B2 => n781, 
                           ZN => n744);
   U1302 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_C_values_1_port, ZN 
                           => n1056);
   U1303 : AOI22D1 port map( A1 => MODE, A2 => n1055, B1 => n1056, B2 => n783, 
                           ZN => n743);
   U1304 : AOI22D1 port map( A1 => MODE, A2 => n1056, B1 => n1057, B2 => n777, 
                           ZN => n742);
   U1305 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_C_values_3_port, ZN 
                           => n1058);
   U1306 : AOI22D1 port map( A1 => MODE, A2 => n1057, B1 => n1058, B2 => n778, 
                           ZN => n741);
   U1307 : AOI22D1 port map( A1 => MODE, A2 => n1058, B1 => n1059, B2 => n782, 
                           ZN => n740);
   U1308 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_C_values_5_port, ZN 
                           => n1060);
   U1309 : AOI22D1 port map( A1 => MODE, A2 => n1059, B1 => n1060, B2 => n782, 
                           ZN => n739);
   U1310 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_C_values_6_port, ZN 
                           => n1061);
   U1311 : AOI22D1 port map( A1 => MODE, A2 => n1060, B1 => n1061, B2 => n782, 
                           ZN => n738);
   U1312 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_C_values_7_port, ZN 
                           => n1062);
   U1313 : AOI22D1 port map( A1 => MODE, A2 => n1061, B1 => n1062, B2 => n782, 
                           ZN => n737);
   U1314 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_C_values_8_port, ZN 
                           => n1063);
   U1315 : AOI22D1 port map( A1 => MODE, A2 => n1062, B1 => n1063, B2 => n782, 
                           ZN => n736);
   U1316 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_C_values_9_port, ZN 
                           => n1064);
   U1317 : AOI22D1 port map( A1 => MODE, A2 => n1063, B1 => n1064, B2 => n782, 
                           ZN => n735);
   U1318 : AOI22D1 port map( A1 => MODE, A2 => n1064, B1 => n1065, B2 => n782, 
                           ZN => n734);
   U1319 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_C_values_11_port, ZN 
                           => n1066);
   U1320 : AOI22D1 port map( A1 => MODE, A2 => n1065, B1 => n1066, B2 => n782, 
                           ZN => n733);
   U1321 : AOI22D1 port map( A1 => MODE, A2 => n1066, B1 => n1067, B2 => n778, 
                           ZN => n732);
   U1322 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_C_values_13_port, ZN 
                           => n1068);
   U1323 : AOI22D1 port map( A1 => MODE, A2 => n1067, B1 => n1068, B2 => n778, 
                           ZN => n731);
   U1324 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_C_values_14_port, ZN 
                           => n1069);
   U1325 : AOI22D1 port map( A1 => MODE, A2 => n1068, B1 => n1069, B2 => n783, 
                           ZN => n730);
   U1326 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_C_values_15_port, ZN 
                           => n1070);
   U1327 : AOI22D1 port map( A1 => MODE, A2 => n1069, B1 => n1070, B2 => n782, 
                           ZN => n729);
   U1328 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_D_values_0_port, ZN 
                           => n1071);
   U1329 : AOI22D1 port map( A1 => MODE, A2 => n1070, B1 => n1071, B2 => n782, 
                           ZN => n728);
   U1330 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_D_values_1_port, ZN 
                           => n1072);
   U1331 : AOI22D1 port map( A1 => MODE, A2 => n1071, B1 => n1072, B2 => n782, 
                           ZN => n727);
   U1332 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_D_values_2_port, ZN 
                           => n1073);
   U1333 : AOI22D1 port map( A1 => MODE, A2 => n1072, B1 => n1073, B2 => n777, 
                           ZN => n726);
   U1334 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_D_values_3_port, ZN 
                           => n1074);
   U1335 : AOI22D1 port map( A1 => MODE, A2 => n1073, B1 => n1074, B2 => n781, 
                           ZN => n725);
   U1336 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_D_values_4_port, ZN 
                           => n1075);
   U1337 : AOI22D1 port map( A1 => MODE, A2 => n1074, B1 => n1075, B2 => n783, 
                           ZN => n724);
   U1338 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_D_values_5_port, ZN 
                           => n1076);
   U1339 : AOI22D1 port map( A1 => MODE, A2 => n1075, B1 => n1076, B2 => n779, 
                           ZN => n723);
   U1340 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_D_values_6_port, ZN 
                           => n1077);
   U1341 : AOI22D1 port map( A1 => MODE, A2 => n1076, B1 => n1077, B2 => n781, 
                           ZN => n722);
   U1342 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_D_values_7_port, ZN 
                           => n1078);
   U1343 : AOI22D1 port map( A1 => MODE, A2 => n1077, B1 => n1078, B2 => n779, 
                           ZN => n721);
   U1344 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_D_values_8_port, ZN 
                           => n1079);
   U1345 : AOI22D1 port map( A1 => MODE, A2 => n1078, B1 => n1079, B2 => n782, 
                           ZN => n720);
   U1346 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_D_values_9_port, ZN 
                           => n1080);
   U1347 : AOI22D1 port map( A1 => MODE, A2 => n1079, B1 => n1080, B2 => n783, 
                           ZN => n719);
   U1348 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_D_values_10_port, ZN 
                           => n1081);
   U1349 : AOI22D1 port map( A1 => MODE, A2 => n1080, B1 => n1081, B2 => n783, 
                           ZN => n718);
   U1350 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_D_values_11_port, ZN 
                           => n1082);
   U1351 : AOI22D1 port map( A1 => MODE, A2 => n1081, B1 => n1082, B2 => n783, 
                           ZN => n717);
   U1352 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_D_values_12_port, ZN 
                           => n1083);
   U1353 : AOI22D1 port map( A1 => MODE, A2 => n1082, B1 => n1083, B2 => n780, 
                           ZN => n716);
   U1354 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_D_values_13_port, ZN 
                           => n1084);
   U1355 : AOI22D1 port map( A1 => MODE, A2 => n1083, B1 => n1084, B2 => n780, 
                           ZN => n715);
   U1356 : INVD0 port map( I => Inst_clb_slice_4xLUT4_LUT_D_values_14_port, ZN 
                           => n1085);
   U1357 : AOI22D1 port map( A1 => MODE, A2 => n1084, B1 => n1085, B2 => n783, 
                           ZN => n714);
   U1358 : INVD0 port map( I => conf_data_1_port, ZN => n1087);
   U1359 : AOI22D1 port map( A1 => MODE, A2 => n1085, B1 => n1087, B2 => n779, 
                           ZN => n713);
   U1360 : AOI22D1 port map( A1 => MODE, A2 => n1087, B1 => n1086, B2 => n783, 
                           ZN => n712);
   U1361 : AOI22D1 port map( A1 => MODE, A2 => n1088, B1 => n524, B2 => n777, 
                           ZN => n709);
   U1362 : AOI22D1 port map( A1 => MODE, A2 => n524, B1 => n527, B2 => n778, ZN
                           => n708);
   U1363 : AOI22D1 port map( A1 => MODE, A2 => n527, B1 => n118, B2 => n780, ZN
                           => n707);
   U1364 : AOI22D1 port map( A1 => MODE, A2 => n118, B1 => n522, B2 => n780, ZN
                           => n706);
   U1365 : AOI22D1 port map( A1 => MODE, A2 => n522, B1 => n1089, B2 => n777, 
                           ZN => n705);
   U1366 : AOI22D1 port map( A1 => MODE, A2 => n1089, B1 => n516, B2 => n778, 
                           ZN => n704);
   U1367 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_173_port, ZN 
                           => n1090);
   U1368 : AOI22D1 port map( A1 => MODE, A2 => n516, B1 => n1090, B2 => n783, 
                           ZN => n703);
   U1369 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_172_port, ZN 
                           => n1091);
   U1370 : AOI22D1 port map( A1 => MODE, A2 => n1090, B1 => n1091, B2 => n778, 
                           ZN => n702);
   U1371 : AOI22D1 port map( A1 => MODE, A2 => n1091, B1 => n127, B2 => n779, 
                           ZN => n701);
   U1372 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_170_port, ZN 
                           => n1092);
   U1373 : AOI22D1 port map( A1 => MODE, A2 => n127, B1 => n1092, B2 => n781, 
                           ZN => n700);
   U1374 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_169_port, ZN 
                           => n1093);
   U1375 : AOI22D1 port map( A1 => MODE, A2 => n1092, B1 => n1093, B2 => n783, 
                           ZN => n699);
   U1376 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_168_port, ZN 
                           => n1094);
   U1377 : AOI22D1 port map( A1 => MODE, A2 => n1093, B1 => n1094, B2 => n779, 
                           ZN => n698);
   U1378 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_167_port, ZN 
                           => n1095);
   U1379 : AOI22D1 port map( A1 => MODE, A2 => n1094, B1 => n1095, B2 => n778, 
                           ZN => n697);
   U1380 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_166_port, ZN 
                           => n1096);
   U1381 : AOI22D1 port map( A1 => MODE, A2 => n1095, B1 => n1096, B2 => n780, 
                           ZN => n696);
   U1382 : AOI22D1 port map( A1 => MODE, A2 => n1096, B1 => n1097, B2 => n780, 
                           ZN => n695);
   U1383 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_164_port, ZN 
                           => n1098);
   U1384 : AOI22D1 port map( A1 => MODE, A2 => n1097, B1 => n1098, B2 => n781, 
                           ZN => n694);
   U1385 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_163_port, ZN 
                           => n1099);
   U1386 : AOI22D1 port map( A1 => MODE, A2 => n1098, B1 => n1099, B2 => n780, 
                           ZN => n693);
   U1387 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_162_port, ZN 
                           => n1100);
   U1388 : AOI22D1 port map( A1 => MODE, A2 => n1099, B1 => n1100, B2 => n780, 
                           ZN => n692);
   U1389 : AOI22D1 port map( A1 => MODE, A2 => n1100, B1 => n136, B2 => n780, 
                           ZN => n691);
   U1390 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_160_port, ZN 
                           => n1101);
   U1391 : AOI22D1 port map( A1 => MODE, A2 => n136, B1 => n1101, B2 => n780, 
                           ZN => n690);
   U1392 : AOI22D1 port map( A1 => MODE, A2 => n1101, B1 => n135, B2 => n780, 
                           ZN => n689);
   U1393 : AOI22D1 port map( A1 => MODE, A2 => n135, B1 => n1102, B2 => n780, 
                           ZN => n688);
   U1394 : AOI22D1 port map( A1 => MODE, A2 => n1102, B1 => n1103, B2 => n780, 
                           ZN => n687);
   U1395 : AOI22D1 port map( A1 => MODE, A2 => n1103, B1 => n505, B2 => n780, 
                           ZN => n686);
   U1396 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_155_port, ZN 
                           => n1104);
   U1397 : AOI22D1 port map( A1 => MODE, A2 => n505, B1 => n1104, B2 => n777, 
                           ZN => n685);
   U1398 : AOI22D1 port map( A1 => MODE, A2 => n1104, B1 => n1105, B2 => n777, 
                           ZN => n684);
   U1399 : AOI22D1 port map( A1 => MODE, A2 => n1105, B1 => n121, B2 => n777, 
                           ZN => n683);
   U1400 : AOI22D1 port map( A1 => MODE, A2 => n121, B1 => n1106, B2 => n777, 
                           ZN => n682);
   U1401 : AOI22D1 port map( A1 => MODE, A2 => n1106, B1 => n1107, B2 => n778, 
                           ZN => n681);
   U1402 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_150_port, ZN 
                           => n1108);
   U1403 : AOI22D1 port map( A1 => MODE, A2 => n1107, B1 => n1108, B2 => n778, 
                           ZN => n680);
   U1404 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_149_port, ZN 
                           => n1109);
   U1405 : AOI22D1 port map( A1 => MODE, A2 => n1108, B1 => n1109, B2 => n777, 
                           ZN => n679);
   U1406 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_148_port, ZN 
                           => n1110);
   U1407 : AOI22D1 port map( A1 => MODE, A2 => n1109, B1 => n1110, B2 => n781, 
                           ZN => n678);
   U1408 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_147_port, ZN 
                           => n1111);
   U1409 : AOI22D1 port map( A1 => MODE, A2 => n1110, B1 => n1111, B2 => n778, 
                           ZN => n677);
   U1410 : AOI22D1 port map( A1 => MODE, A2 => n1111, B1 => n1112, B2 => n777, 
                           ZN => n676);
   U1411 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_145_port, ZN 
                           => n1113);
   U1412 : AOI22D1 port map( A1 => MODE, A2 => n1112, B1 => n1113, B2 => n777, 
                           ZN => n675);
   U1413 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_144_port, ZN 
                           => n1114);
   U1414 : AOI22D1 port map( A1 => MODE, A2 => n1113, B1 => n1114, B2 => n782, 
                           ZN => n674);
   U1415 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_143_port, ZN 
                           => n1115);
   U1416 : AOI22D1 port map( A1 => MODE, A2 => n1114, B1 => n1115, B2 => n777, 
                           ZN => n673);
   U1417 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_142_port, ZN 
                           => n1116);
   U1418 : AOI22D1 port map( A1 => MODE, A2 => n1115, B1 => n1116, B2 => n779, 
                           ZN => n672);
   U1419 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_141_port, ZN 
                           => n1117);
   U1420 : AOI22D1 port map( A1 => MODE, A2 => n1116, B1 => n1117, B2 => n780, 
                           ZN => n671);
   U1421 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_140_port, ZN 
                           => n1118);
   U1422 : AOI22D1 port map( A1 => MODE, A2 => n1117, B1 => n1118, B2 => n777, 
                           ZN => n670);
   U1423 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_139_port, ZN 
                           => n1119);
   U1424 : AOI22D1 port map( A1 => MODE, A2 => n1118, B1 => n1119, B2 => n778, 
                           ZN => n669);
   U1425 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_138_port, ZN 
                           => n1120);
   U1426 : AOI22D1 port map( A1 => MODE, A2 => n1119, B1 => n1120, B2 => n781, 
                           ZN => n668);
   U1427 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_137_port, ZN 
                           => n1121);
   U1428 : AOI22D1 port map( A1 => MODE, A2 => n1120, B1 => n1121, B2 => n778, 
                           ZN => n667);
   U1429 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_136_port, ZN 
                           => n1122);
   U1430 : AOI22D1 port map( A1 => MODE, A2 => n1121, B1 => n1122, B2 => n778, 
                           ZN => n666);
   U1431 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_135_port, ZN 
                           => n1123);
   U1432 : AOI22D1 port map( A1 => MODE, A2 => n1122, B1 => n1123, B2 => n778, 
                           ZN => n665);
   U1433 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_134_port, ZN 
                           => n1124);
   U1434 : AOI22D1 port map( A1 => MODE, A2 => n1123, B1 => n1124, B2 => n778, 
                           ZN => n664);
   U1435 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_133_port, ZN 
                           => n1125);
   U1436 : AOI22D1 port map( A1 => MODE, A2 => n1124, B1 => n1125, B2 => n778, 
                           ZN => n663);
   U1437 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_132_port, ZN 
                           => n1126);
   U1438 : AOI22D1 port map( A1 => MODE, A2 => n1125, B1 => n1126, B2 => n778, 
                           ZN => n662);
   U1439 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_131_port, ZN 
                           => n1127);
   U1440 : AOI22D1 port map( A1 => MODE, A2 => n1126, B1 => n1127, B2 => n777, 
                           ZN => n661);
   U1441 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_130_port, ZN 
                           => n1128);
   U1442 : AOI22D1 port map( A1 => MODE, A2 => n1127, B1 => n1128, B2 => n778, 
                           ZN => n660);
   U1443 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_129_port, ZN 
                           => n1129);
   U1444 : AOI22D1 port map( A1 => MODE, A2 => n1128, B1 => n1129, B2 => n777, 
                           ZN => n659);
   U1445 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_128_port, ZN 
                           => n1130);
   U1446 : AOI22D1 port map( A1 => MODE, A2 => n1129, B1 => n1130, B2 => n778, 
                           ZN => n658);
   U1447 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_127_port, ZN 
                           => n1131);
   U1448 : AOI22D1 port map( A1 => MODE, A2 => n1130, B1 => n1131, B2 => n783, 
                           ZN => n657);
   U1449 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_126_port, ZN 
                           => n1132);
   U1450 : AOI22D1 port map( A1 => MODE, A2 => n1131, B1 => n1132, B2 => n779, 
                           ZN => n656);
   U1451 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_125_port, ZN 
                           => n1133);
   U1452 : AOI22D1 port map( A1 => MODE, A2 => n1132, B1 => n1133, B2 => n778, 
                           ZN => n655);
   U1453 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_124_port, ZN 
                           => n1134);
   U1454 : AOI22D1 port map( A1 => MODE, A2 => n1133, B1 => n1134, B2 => n781, 
                           ZN => n654);
   U1455 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_123_port, ZN 
                           => n1135);
   U1456 : AOI22D1 port map( A1 => MODE, A2 => n1134, B1 => n1135, B2 => n781, 
                           ZN => n653);
   U1457 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_122_port, ZN 
                           => n1136);
   U1458 : AOI22D1 port map( A1 => MODE, A2 => n1135, B1 => n1136, B2 => n780, 
                           ZN => n652);
   U1459 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_121_port, ZN 
                           => n1137);
   U1460 : AOI22D1 port map( A1 => MODE, A2 => n1136, B1 => n1137, B2 => n779, 
                           ZN => n651);
   U1461 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_120_port, ZN 
                           => n1138);
   U1462 : AOI22D1 port map( A1 => MODE, A2 => n1137, B1 => n1138, B2 => n777, 
                           ZN => n650);
   U1463 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_119_port, ZN 
                           => n1139);
   U1464 : AOI22D1 port map( A1 => MODE, A2 => n1138, B1 => n1139, B2 => n778, 
                           ZN => n649);
   U1465 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_118_port, ZN 
                           => n1140);
   U1466 : AOI22D1 port map( A1 => MODE, A2 => n1139, B1 => n1140, B2 => n777, 
                           ZN => n648);
   U1467 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_117_port, ZN 
                           => n1141);
   U1468 : AOI22D1 port map( A1 => MODE, A2 => n1140, B1 => n1141, B2 => n778, 
                           ZN => n647);
   U1469 : AOI22D1 port map( A1 => MODE, A2 => n1141, B1 => n1142, B2 => n783, 
                           ZN => n646);
   U1470 : AOI22D1 port map( A1 => MODE, A2 => n1142, B1 => n1143, B2 => n780, 
                           ZN => n645);
   U1471 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_114_port, ZN 
                           => n1144);
   U1472 : AOI22D1 port map( A1 => MODE, A2 => n1143, B1 => n1144, B2 => n778, 
                           ZN => n644);
   U1473 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_113_port, ZN 
                           => n1145);
   U1474 : AOI22D1 port map( A1 => MODE, A2 => n1144, B1 => n1145, B2 => n777, 
                           ZN => n643);
   U1475 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_112_port, ZN 
                           => n1146);
   U1476 : AOI22D1 port map( A1 => MODE, A2 => n1145, B1 => n1146, B2 => n783, 
                           ZN => n642);
   U1477 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_111_port, ZN 
                           => n1147);
   U1478 : AOI22D1 port map( A1 => MODE, A2 => n1146, B1 => n1147, B2 => n781, 
                           ZN => n641);
   U1479 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_110_port, ZN 
                           => n1148);
   U1480 : AOI22D1 port map( A1 => MODE, A2 => n1147, B1 => n1148, B2 => n782, 
                           ZN => n640);
   U1481 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_109_port, ZN 
                           => n1149);
   U1482 : AOI22D1 port map( A1 => MODE, A2 => n1148, B1 => n1149, B2 => n777, 
                           ZN => n639);
   U1483 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_108_port, ZN 
                           => n1150);
   U1484 : AOI22D1 port map( A1 => MODE, A2 => n1149, B1 => n1150, B2 => n780, 
                           ZN => n638);
   U1485 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_107_port, ZN 
                           => n1151);
   U1486 : AOI22D1 port map( A1 => MODE, A2 => n1150, B1 => n1151, B2 => n778, 
                           ZN => n637);
   U1487 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_106_port, ZN 
                           => n1152);
   U1488 : AOI22D1 port map( A1 => MODE, A2 => n1151, B1 => n1152, B2 => n779, 
                           ZN => n636);
   U1489 : AOI22D1 port map( A1 => MODE, A2 => n1152, B1 => n1153, B2 => n782, 
                           ZN => n635);
   U1490 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_104_port, ZN 
                           => n1154);
   U1491 : AOI22D1 port map( A1 => MODE, A2 => n1153, B1 => n1154, B2 => n783, 
                           ZN => n634);
   U1492 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_103_port, ZN 
                           => n1155);
   U1493 : AOI22D1 port map( A1 => MODE, A2 => n1154, B1 => n1155, B2 => n783, 
                           ZN => n633);
   U1494 : AOI22D1 port map( A1 => MODE, A2 => n1155, B1 => n1156, B2 => n777, 
                           ZN => n632);
   U1495 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_101_port, ZN 
                           => n1157);
   U1496 : AOI22D1 port map( A1 => MODE, A2 => n1156, B1 => n1157, B2 => n783, 
                           ZN => n631);
   U1497 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_100_port, ZN 
                           => n1158);
   U1498 : AOI22D1 port map( A1 => MODE, A2 => n1157, B1 => n1158, B2 => n778, 
                           ZN => n630);
   U1499 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_99_port, ZN 
                           => n1159);
   U1500 : AOI22D1 port map( A1 => MODE, A2 => n1158, B1 => n1159, B2 => n779, 
                           ZN => n629);
   U1501 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_98_port, ZN 
                           => n1160);
   U1502 : AOI22D1 port map( A1 => MODE, A2 => n1159, B1 => n1160, B2 => n782, 
                           ZN => n628);
   U1503 : AOI22D1 port map( A1 => MODE, A2 => n1160, B1 => n1161, B2 => n783, 
                           ZN => n627);
   U1504 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_96_port, ZN 
                           => n1162);
   U1505 : AOI22D1 port map( A1 => MODE, A2 => n1161, B1 => n1162, B2 => n783, 
                           ZN => n626);
   U1506 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_95_port, ZN 
                           => n1163);
   U1507 : AOI22D1 port map( A1 => MODE, A2 => n1162, B1 => n1163, B2 => n781, 
                           ZN => n625);
   U1508 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_94_port, ZN 
                           => n1164);
   U1509 : AOI22D1 port map( A1 => MODE, A2 => n1163, B1 => n1164, B2 => n781, 
                           ZN => n624);
   U1510 : AOI22D1 port map( A1 => MODE, A2 => n1164, B1 => n1165, B2 => n782, 
                           ZN => n623);
   U1511 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_92_port, ZN 
                           => n1166);
   U1512 : AOI22D1 port map( A1 => MODE, A2 => n1165, B1 => n1166, B2 => n778, 
                           ZN => n622);
   U1513 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_91_port, ZN 
                           => n1167);
   U1514 : AOI22D1 port map( A1 => MODE, A2 => n1166, B1 => n1167, B2 => n781, 
                           ZN => n621);
   U1515 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_90_port, ZN 
                           => n1168);
   U1516 : AOI22D1 port map( A1 => MODE, A2 => n1167, B1 => n1168, B2 => n779, 
                           ZN => n620);
   U1517 : AOI22D1 port map( A1 => MODE, A2 => n1168, B1 => n1169, B2 => n778, 
                           ZN => n619);
   U1518 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_88_port, ZN 
                           => n1170);
   U1519 : AOI22D1 port map( A1 => MODE, A2 => n1169, B1 => n1170, B2 => n779, 
                           ZN => n618);
   U1520 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_87_port, ZN 
                           => n1171);
   U1521 : AOI22D1 port map( A1 => MODE, A2 => n1170, B1 => n1171, B2 => n778, 
                           ZN => n617);
   U1522 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_86_port, ZN 
                           => n1172);
   U1523 : AOI22D1 port map( A1 => MODE, A2 => n1171, B1 => n1172, B2 => n783, 
                           ZN => n616);
   U1524 : AOI22D1 port map( A1 => MODE, A2 => n1172, B1 => n1173, B2 => n777, 
                           ZN => n615);
   U1525 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_84_port, ZN 
                           => n1174);
   U1526 : AOI22D1 port map( A1 => MODE, A2 => n1173, B1 => n1174, B2 => n783, 
                           ZN => n614);
   U1527 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_83_port, ZN 
                           => n1175);
   U1528 : AOI22D1 port map( A1 => MODE, A2 => n1174, B1 => n1175, B2 => n777, 
                           ZN => n613);
   U1529 : AOI22D1 port map( A1 => MODE, A2 => n1175, B1 => n1176, B2 => n783, 
                           ZN => n612);
   U1530 : AOI22D1 port map( A1 => MODE, A2 => n1176, B1 => n1177, B2 => n778, 
                           ZN => n611);
   U1531 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_80_port, ZN 
                           => n1178);
   U1532 : AOI22D1 port map( A1 => MODE, A2 => n1177, B1 => n1178, B2 => n780, 
                           ZN => n610);
   U1533 : AOI22D1 port map( A1 => MODE, A2 => n1178, B1 => n1179, B2 => n782, 
                           ZN => n609);
   U1534 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_78_port, ZN 
                           => n1180);
   U1535 : AOI22D1 port map( A1 => MODE, A2 => n1179, B1 => n1180, B2 => n778, 
                           ZN => n608);
   U1536 : AOI22D1 port map( A1 => MODE, A2 => n1180, B1 => n1181, B2 => n777, 
                           ZN => n607);
   U1537 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_76_port, ZN 
                           => n1182);
   U1538 : AOI22D1 port map( A1 => MODE, A2 => n1181, B1 => n1182, B2 => n778, 
                           ZN => n606);
   U1539 : AOI22D1 port map( A1 => MODE, A2 => n1182, B1 => n1183, B2 => n781, 
                           ZN => n605);
   U1540 : AOI22D1 port map( A1 => MODE, A2 => n1183, B1 => n1184, B2 => n779, 
                           ZN => n604);
   U1541 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_73_port, ZN 
                           => n1185);
   U1542 : AOI22D1 port map( A1 => MODE, A2 => n1184, B1 => n1185, B2 => n781, 
                           ZN => n603);
   U1543 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_72_port, ZN 
                           => n1186);
   U1544 : AOI22D1 port map( A1 => MODE, A2 => n1185, B1 => n1186, B2 => n783, 
                           ZN => n602);
   U1545 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_71_port, ZN 
                           => n1187);
   U1546 : AOI22D1 port map( A1 => MODE, A2 => n1186, B1 => n1187, B2 => n777, 
                           ZN => n601);
   U1547 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_70_port, ZN 
                           => n1188);
   U1548 : AOI22D1 port map( A1 => MODE, A2 => n1187, B1 => n1188, B2 => n779, 
                           ZN => n600);
   U1549 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_69_port, ZN 
                           => n1189);
   U1550 : AOI22D1 port map( A1 => MODE, A2 => n1188, B1 => n1189, B2 => n781, 
                           ZN => n599);
   U1551 : AOI22D1 port map( A1 => MODE, A2 => n1189, B1 => n1190, B2 => n778, 
                           ZN => n598);
   U1552 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_67_port, ZN 
                           => n1191);
   U1553 : AOI22D1 port map( A1 => MODE, A2 => n1190, B1 => n1191, B2 => n779, 
                           ZN => n597);
   U1554 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_66_port, ZN 
                           => n1192);
   U1555 : AOI22D1 port map( A1 => MODE, A2 => n1191, B1 => n1192, B2 => n781, 
                           ZN => n596);
   U1556 : AOI22D1 port map( A1 => MODE, A2 => n1192, B1 => n1193, B2 => n779, 
                           ZN => n595);
   U1557 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_64_port, ZN 
                           => n1194);
   U1558 : AOI22D1 port map( A1 => MODE, A2 => n1193, B1 => n1194, B2 => n781, 
                           ZN => n594);
   U1559 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_63_port, ZN 
                           => n1195);
   U1560 : AOI22D1 port map( A1 => MODE, A2 => n1194, B1 => n1195, B2 => n783, 
                           ZN => n593);
   U1561 : AOI22D1 port map( A1 => MODE, A2 => n1195, B1 => n1196, B2 => n778, 
                           ZN => n592);
   U1562 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_61_port, ZN 
                           => n1197);
   U1563 : AOI22D1 port map( A1 => MODE, A2 => n1196, B1 => n1197, B2 => n777, 
                           ZN => n591);
   U1564 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_60_port, ZN 
                           => n1198);
   U1565 : AOI22D1 port map( A1 => MODE, A2 => n1197, B1 => n1198, B2 => n778, 
                           ZN => n590);
   U1566 : AOI22D1 port map( A1 => MODE, A2 => n1198, B1 => n1199, B2 => n777, 
                           ZN => n589);
   U1567 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_58_port, ZN 
                           => n1200);
   U1568 : AOI22D1 port map( A1 => MODE, A2 => n1199, B1 => n1200, B2 => n777, 
                           ZN => n588);
   U1569 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_57_port, ZN 
                           => n1201);
   U1570 : AOI22D1 port map( A1 => MODE, A2 => n1200, B1 => n1201, B2 => n777, 
                           ZN => n587);
   U1571 : AOI22D1 port map( A1 => MODE, A2 => n1201, B1 => n1202, B2 => n778, 
                           ZN => n586);
   U1572 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_55_port, ZN 
                           => n1203);
   U1573 : AOI22D1 port map( A1 => MODE, A2 => n1202, B1 => n1203, B2 => n777, 
                           ZN => n585);
   U1574 : AOI22D1 port map( A1 => MODE, A2 => n1203, B1 => n1204, B2 => n783, 
                           ZN => n584);
   U1575 : AOI22D1 port map( A1 => MODE, A2 => n1204, B1 => n1205, B2 => n782, 
                           ZN => n583);
   U1576 : AOI22D1 port map( A1 => MODE, A2 => n1205, B1 => n1206, B2 => n777, 
                           ZN => n582);
   U1577 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_51_port, ZN 
                           => n1207);
   U1578 : AOI22D1 port map( A1 => MODE, A2 => n1206, B1 => n1207, B2 => n783, 
                           ZN => n581);
   U1579 : AOI22D1 port map( A1 => MODE, A2 => n1207, B1 => n1208, B2 => n777, 
                           ZN => n580);
   U1580 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_49_port, ZN 
                           => n1209);
   U1581 : AOI22D1 port map( A1 => MODE, A2 => n1208, B1 => n1209, B2 => n777, 
                           ZN => n579);
   U1582 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_48_port, ZN 
                           => n1210);
   U1583 : AOI22D1 port map( A1 => MODE, A2 => n1209, B1 => n1210, B2 => n777, 
                           ZN => n578);
   U1584 : AOI22D1 port map( A1 => MODE, A2 => n1210, B1 => n1211, B2 => n780, 
                           ZN => n577);
   U1585 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_46_port, ZN 
                           => n1212);
   U1586 : AOI22D1 port map( A1 => MODE, A2 => n1211, B1 => n1212, B2 => n779, 
                           ZN => n576);
   U1587 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_45_port, ZN 
                           => n1213);
   U1588 : AOI22D1 port map( A1 => MODE, A2 => n1212, B1 => n1213, B2 => n781, 
                           ZN => n575);
   U1589 : AOI22D1 port map( A1 => MODE, A2 => n1213, B1 => n1214, B2 => n778, 
                           ZN => n574);
   U1590 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_43_port, ZN 
                           => n1215);
   U1591 : AOI22D1 port map( A1 => MODE, A2 => n1214, B1 => n1215, B2 => n782, 
                           ZN => n573);
   U1592 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_42_port, ZN 
                           => n1216);
   U1593 : AOI22D1 port map( A1 => MODE, A2 => n1215, B1 => n1216, B2 => n777, 
                           ZN => n572);
   U1594 : AOI22D1 port map( A1 => MODE, A2 => n1216, B1 => n1217, B2 => n778, 
                           ZN => n571);
   U1595 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_40_port, ZN 
                           => n1218);
   U1596 : AOI22D1 port map( A1 => MODE, A2 => n1217, B1 => n1218, B2 => n777, 
                           ZN => n570);
   U1597 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_39_port, ZN 
                           => n1219);
   U1598 : AOI22D1 port map( A1 => MODE, A2 => n1218, B1 => n1219, B2 => n778, 
                           ZN => n569);
   U1599 : AOI22D1 port map( A1 => MODE, A2 => n1219, B1 => n1220, B2 => n778, 
                           ZN => n568);
   U1600 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_37_port, ZN 
                           => n1221);
   U1601 : AOI22D1 port map( A1 => MODE, A2 => n1220, B1 => n1221, B2 => n781, 
                           ZN => n567);
   U1602 : AOI22D1 port map( A1 => MODE, A2 => n1221, B1 => n1222, B2 => n777, 
                           ZN => n566);
   U1603 : AOI22D1 port map( A1 => MODE, A2 => n1222, B1 => n1223, B2 => n777, 
                           ZN => n565);
   U1604 : AOI22D1 port map( A1 => MODE, A2 => n1223, B1 => n1224, B2 => n777, 
                           ZN => n564);
   U1605 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_33_port, ZN 
                           => n1225);
   U1606 : AOI22D1 port map( A1 => MODE, A2 => n1224, B1 => n1225, B2 => n780, 
                           ZN => n563);
   U1607 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_32_port, ZN 
                           => n1226);
   U1608 : AOI22D1 port map( A1 => MODE, A2 => n1225, B1 => n1226, B2 => n777, 
                           ZN => n562);
   U1609 : AOI22D1 port map( A1 => MODE, A2 => n1226, B1 => n1227, B2 => n779, 
                           ZN => n561);
   U1610 : AOI22D1 port map( A1 => MODE, A2 => n1227, B1 => n1228, B2 => n779, 
                           ZN => n560);
   U1611 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_29_port, ZN 
                           => n1229);
   U1612 : AOI22D1 port map( A1 => MODE, A2 => n1228, B1 => n1229, B2 => n777, 
                           ZN => n559);
   U1613 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_28_port, ZN 
                           => n1230);
   U1614 : AOI22D1 port map( A1 => MODE, A2 => n1229, B1 => n1230, B2 => n778, 
                           ZN => n558);
   U1615 : AOI22D1 port map( A1 => MODE, A2 => n1230, B1 => n1231, B2 => n783, 
                           ZN => n557);
   U1616 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_26_port, ZN 
                           => n1232);
   U1617 : AOI22D1 port map( A1 => MODE, A2 => n1231, B1 => n1232, B2 => n781, 
                           ZN => n556);
   U1618 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_25_port, ZN 
                           => n1233);
   U1619 : AOI22D1 port map( A1 => MODE, A2 => n1232, B1 => n1233, B2 => n782, 
                           ZN => n555);
   U1620 : AOI22D1 port map( A1 => MODE, A2 => n1233, B1 => n1234, B2 => n782, 
                           ZN => n554);
   U1621 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_23_port, ZN 
                           => n1235);
   U1622 : AOI22D1 port map( A1 => MODE, A2 => n1234, B1 => n1235, B2 => n782, 
                           ZN => n553);
   U1623 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_22_port, ZN 
                           => n1236);
   U1624 : AOI22D1 port map( A1 => MODE, A2 => n1235, B1 => n1236, B2 => n779, 
                           ZN => n552);
   U1625 : AOI22D1 port map( A1 => MODE, A2 => n1236, B1 => n1237, B2 => n781, 
                           ZN => n551);
   U1626 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_20_port, ZN 
                           => n1238);
   U1627 : AOI22D1 port map( A1 => MODE, A2 => n1237, B1 => n1238, B2 => n779, 
                           ZN => n550);
   U1628 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_19_port, ZN 
                           => n1239);
   U1629 : AOI22D1 port map( A1 => MODE, A2 => n1238, B1 => n1239, B2 => n783, 
                           ZN => n549);
   U1630 : AOI22D1 port map( A1 => MODE, A2 => n1239, B1 => n1240, B2 => n777, 
                           ZN => n548);
   U1631 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_17_port, ZN 
                           => n1241);
   U1632 : AOI22D1 port map( A1 => MODE, A2 => n1240, B1 => n1241, B2 => n778, 
                           ZN => n547);
   U1633 : AOI22D1 port map( A1 => MODE, A2 => n1241, B1 => n1242, B2 => n778, 
                           ZN => n546);
   U1634 : AOI22D1 port map( A1 => MODE, A2 => n1242, B1 => n1243, B2 => n777, 
                           ZN => n545);
   U1635 : AOI22D1 port map( A1 => MODE, A2 => n1243, B1 => n1244, B2 => n777, 
                           ZN => n544);
   U1636 : AOI22D1 port map( A1 => MODE, A2 => n1244, B1 => n1245, B2 => n781, 
                           ZN => n543);
   U1637 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_12_port, ZN 
                           => n1246);
   U1638 : AOI22D1 port map( A1 => MODE, A2 => n1245, B1 => n1246, B2 => n779, 
                           ZN => n542);
   U1639 : AOI22D1 port map( A1 => MODE, A2 => n1246, B1 => n1247, B2 => n782, 
                           ZN => n541);
   U1640 : AOI22D1 port map( A1 => MODE, A2 => n1247, B1 => n1248, B2 => n778, 
                           ZN => n540);
   U1641 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_9_port, ZN =>
                           n1249);
   U1642 : AOI22D1 port map( A1 => MODE, A2 => n1248, B1 => n1249, B2 => n780, 
                           ZN => n539);
   U1643 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_8_port, ZN =>
                           n1250);
   U1644 : AOI22D1 port map( A1 => MODE, A2 => n1249, B1 => n1250, B2 => n779, 
                           ZN => n538);
   U1645 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_7_port, ZN =>
                           n1251);
   U1646 : AOI22D1 port map( A1 => MODE, A2 => n1250, B1 => n1251, B2 => n781, 
                           ZN => n537);
   U1647 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_6_port, ZN =>
                           n1252);
   U1648 : AOI22D1 port map( A1 => MODE, A2 => n1251, B1 => n1252, B2 => n779, 
                           ZN => n536);
   U1649 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_5_port, ZN =>
                           n1253);
   U1650 : AOI22D1 port map( A1 => MODE, A2 => n1252, B1 => n1253, B2 => n780, 
                           ZN => n535);
   U1651 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_4_port, ZN =>
                           n1254);
   U1652 : AOI22D1 port map( A1 => MODE, A2 => n1253, B1 => n1254, B2 => n779, 
                           ZN => n534);
   U1653 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_3_port, ZN =>
                           n1255);
   U1654 : AOI22D1 port map( A1 => MODE, A2 => n1254, B1 => n1255, B2 => n779, 
                           ZN => n533);
   U1655 : INVD0 port map( I => Inst_CLB_switch_matrix_ConfigBits_2_port, ZN =>
                           n1257);
   U1656 : AOI22D1 port map( A1 => MODE, A2 => n1255, B1 => n1257, B2 => n778, 
                           ZN => n532);
   U1657 : AOI22D1 port map( A1 => MODE, A2 => n1257, B1 => n1256, B2 => n781, 
                           ZN => n531);
   U1658 : MUX4D1 port map( I0 => IJ_BEG_8_port, I1 => IJ_BEG_10_port, I2 => 
                           IJ_BEG_9_port, I3 => IJ_BEG_11_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_148_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_147_port, Z => 
                           IJ_BEG_0_port);
   U1659 : MUX4D1 port map( I0 => IJ_BEG_6_port, I1 => IJ_BEG_8_port, I2 => 
                           IJ_BEG_7_port, I3 => IJ_BEG_9_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_144_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_143_port, Z => D3)
                           ;
   U1660 : MUX4D1 port map( I0 => IJ_BEG_5_port, I1 => IJ_BEG_7_port, I2 => 
                           IJ_BEG_6_port, I3 => IJ_BEG_8_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_142_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_141_port, Z => D2)
                           ;
   U1661 : MUX4D1 port map( I0 => IJ_BEG_4_port, I1 => IJ_BEG_6_port, I2 => 
                           IJ_BEG_5_port, I3 => IJ_BEG_7_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_140_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_139_port, Z => D1)
                           ;
   U1662 : MUX4D1 port map( I0 => IJ_BEG_3_port, I1 => IJ_BEG_5_port, I2 => 
                           IJ_BEG_4_port, I3 => IJ_BEG_6_port, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_138_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_137_port, Z => D0)
                           ;
   U1663 : MUX4D1 port map( I0 => A, I1 => B, I2 => AQ, I3 => BQ, S0 => 
                           Inst_CLB_switch_matrix_ConfigBits_114_port, S1 => 
                           Inst_CLB_switch_matrix_ConfigBits_113_port, Z => A0)
                           ;

end SYN_Behavioral;
