//NumberOfConfigBits:406
module DSP_top_switch_matrix (N1END0, N1END1, N1END2, N1END3, N2MID0, N2MID1, N2MID2, N2MID3, N2MID4, N2MID5, N2MID6, N2MID7, N2END0, N2END1, N2END2, N2END3, N2END4, N2END5, N2END6, N2END7, N4END0, N4END1, N4END2, N4END3, NN4END0, NN4END1, NN4END2, NN4END3, bot2top0, bot2top1, bot2top2, bot2top3, bot2top4, bot2top5, bot2top6, bot2top7, bot2top8, bot2top9, E1END0, E1END1, E1END2, E1END3, E2MID0, E2MID1, E2MID2, E2MID3, E2MID4, E2MID5, E2MID6, E2MID7, E2END0, E2END1, E2END2, E2END3, E2END4, E2END5, E2END6, E2END7, EE4END0, EE4END1, EE4END2, EE4END3, E6END0, E6END1, S1END0, S1END1, S1END2, S1END3, S2MID0, S2MID1, S2MID2, S2MID3, S2MID4, S2MID5, S2MID6, S2MID7, S2END0, S2END1, S2END2, S2END3, S2END4, S2END5, S2END6, S2END7, S4END0, S4END1, S4END2, S4END3, SS4END0, SS4END1, SS4END2, SS4END3, W1END0, W1END1, W1END2, W1END3, W2MID0, W2MID1, W2MID2, W2MID3, W2MID4, W2MID5, W2MID6, W2MID7, W2END0, W2END1, W2END2, W2END3, W2END4, W2END5, W2END6, W2END7, WW4END0, WW4END1, WW4END2, WW4END3, W6END0, W6END1, J2MID_ABa_END0, J2MID_ABa_END1, J2MID_ABa_END2, J2MID_ABa_END3, J2MID_CDa_END0, J2MID_CDa_END1, J2MID_CDa_END2, J2MID_CDa_END3, J2MID_EFa_END0, J2MID_EFa_END1, J2MID_EFa_END2, J2MID_EFa_END3, J2MID_GHa_END0, J2MID_GHa_END1, J2MID_GHa_END2, J2MID_GHa_END3, J2MID_ABb_END0, J2MID_ABb_END1, J2MID_ABb_END2, J2MID_ABb_END3, J2MID_CDb_END0, J2MID_CDb_END1, J2MID_CDb_END2, J2MID_CDb_END3, J2MID_EFb_END0, J2MID_EFb_END1, J2MID_EFb_END2, J2MID_EFb_END3, J2MID_GHb_END0, J2MID_GHb_END1, J2MID_GHb_END2, J2MID_GHb_END3, J2END_AB_END0, J2END_AB_END1, J2END_AB_END2, J2END_AB_END3, J2END_CD_END0, J2END_CD_END1, J2END_CD_END2, J2END_CD_END3, J2END_EF_END0, J2END_EF_END1, J2END_EF_END2, J2END_EF_END3, J2END_GH_END0, J2END_GH_END1, J2END_GH_END2, J2END_GH_END3, JN2END0, JN2END1, JN2END2, JN2END3, JN2END4, JN2END5, JN2END6, JN2END7, JE2END0, JE2END1, JE2END2, JE2END3, JE2END4, JE2END5, JE2END6, JE2END7, JS2END0, JS2END1, JS2END2, JS2END3, JS2END4, JS2END5, JS2END6, JS2END7, JW2END0, JW2END1, JW2END2, JW2END3, JW2END4, JW2END5, JW2END6, JW2END7, J_l_AB_END0, J_l_AB_END1, J_l_AB_END2, J_l_AB_END3, J_l_CD_END0, J_l_CD_END1, J_l_CD_END2, J_l_CD_END3, J_l_EF_END0, J_l_EF_END1, J_l_EF_END2, J_l_EF_END3, J_l_GH_END0, J_l_GH_END1, J_l_GH_END2, J_l_GH_END3, N1BEG0, N1BEG1, N1BEG2, N1BEG3, N2BEG0, N2BEG1, N2BEG2, N2BEG3, N2BEG4, N2BEG5, N2BEG6, N2BEG7, N2BEGb0, N2BEGb1, N2BEGb2, N2BEGb3, N2BEGb4, N2BEGb5, N2BEGb6, N2BEGb7, N4BEG0, N4BEG1, N4BEG2, N4BEG3, NN4BEG0, NN4BEG1, NN4BEG2, NN4BEG3, E1BEG0, E1BEG1, E1BEG2, E1BEG3, E2BEG0, E2BEG1, E2BEG2, E2BEG3, E2BEG4, E2BEG5, E2BEG6, E2BEG7, E2BEGb0, E2BEGb1, E2BEGb2, E2BEGb3, E2BEGb4, E2BEGb5, E2BEGb6, E2BEGb7, EE4BEG0, EE4BEG1, EE4BEG2, EE4BEG3, E6BEG0, E6BEG1, S1BEG0, S1BEG1, S1BEG2, S1BEG3, S2BEG0, S2BEG1, S2BEG2, S2BEG3, S2BEG4, S2BEG5, S2BEG6, S2BEG7, S2BEGb0, S2BEGb1, S2BEGb2, S2BEGb3, S2BEGb4, S2BEGb5, S2BEGb6, S2BEGb7, S4BEG0, S4BEG1, S4BEG2, S4BEG3, SS4BEG0, SS4BEG1, SS4BEG2, SS4BEG3, top2bot0, top2bot1, top2bot2, top2bot3, top2bot4, top2bot5, top2bot6, top2bot7, top2bot8, top2bot9, top2bot10, top2bot11, top2bot12, top2bot13, top2bot14, top2bot15, top2bot16, top2bot17, W1BEG0, W1BEG1, W1BEG2, W1BEG3, W2BEG0, W2BEG1, W2BEG2, W2BEG3, W2BEG4, W2BEG5, W2BEG6, W2BEG7, W2BEGb0, W2BEGb1, W2BEGb2, W2BEGb3, W2BEGb4, W2BEGb5, W2BEGb6, W2BEGb7, WW4BEG0, WW4BEG1, WW4BEG2, WW4BEG3, W6BEG0, W6BEG1, J2MID_ABa_BEG0, J2MID_ABa_BEG1, J2MID_ABa_BEG2, J2MID_ABa_BEG3, J2MID_CDa_BEG0, J2MID_CDa_BEG1, J2MID_CDa_BEG2, J2MID_CDa_BEG3, J2MID_EFa_BEG0, J2MID_EFa_BEG1, J2MID_EFa_BEG2, J2MID_EFa_BEG3, J2MID_GHa_BEG0, J2MID_GHa_BEG1, J2MID_GHa_BEG2, J2MID_GHa_BEG3, J2MID_ABb_BEG0, J2MID_ABb_BEG1, J2MID_ABb_BEG2, J2MID_ABb_BEG3, J2MID_CDb_BEG0, J2MID_CDb_BEG1, J2MID_CDb_BEG2, J2MID_CDb_BEG3, J2MID_EFb_BEG0, J2MID_EFb_BEG1, J2MID_EFb_BEG2, J2MID_EFb_BEG3, J2MID_GHb_BEG0, J2MID_GHb_BEG1, J2MID_GHb_BEG2, J2MID_GHb_BEG3, J2END_AB_BEG0, J2END_AB_BEG1, J2END_AB_BEG2, J2END_AB_BEG3, J2END_CD_BEG0, J2END_CD_BEG1, J2END_CD_BEG2, J2END_CD_BEG3, J2END_EF_BEG0, J2END_EF_BEG1, J2END_EF_BEG2, J2END_EF_BEG3, J2END_GH_BEG0, J2END_GH_BEG1, J2END_GH_BEG2, J2END_GH_BEG3, JN2BEG0, JN2BEG1, JN2BEG2, JN2BEG3, JN2BEG4, JN2BEG5, JN2BEG6, JN2BEG7, JE2BEG0, JE2BEG1, JE2BEG2, JE2BEG3, JE2BEG4, JE2BEG5, JE2BEG6, JE2BEG7, JS2BEG0, JS2BEG1, JS2BEG2, JS2BEG3, JS2BEG4, JS2BEG5, JS2BEG6, JS2BEG7, JW2BEG0, JW2BEG1, JW2BEG2, JW2BEG3, JW2BEG4, JW2BEG5, JW2BEG6, JW2BEG7, J_l_AB_BEG0, J_l_AB_BEG1, J_l_AB_BEG2, J_l_AB_BEG3, J_l_CD_BEG0, J_l_CD_BEG1, J_l_CD_BEG2, J_l_CD_BEG3, J_l_EF_BEG0, J_l_EF_BEG1, J_l_EF_BEG2, J_l_EF_BEG3, J_l_GH_BEG0, J_l_GH_BEG1, J_l_GH_BEG2, J_l_GH_BEG3, ConfigBits, ConfigBits_N);
	parameter NoConfigBits = 406;
	 // switch matrix inputs
	input N1END0;
	input N1END1;
	input N1END2;
	input N1END3;
	input N2MID0;
	input N2MID1;
	input N2MID2;
	input N2MID3;
	input N2MID4;
	input N2MID5;
	input N2MID6;
	input N2MID7;
	input N2END0;
	input N2END1;
	input N2END2;
	input N2END3;
	input N2END4;
	input N2END5;
	input N2END6;
	input N2END7;
	input N4END0;
	input N4END1;
	input N4END2;
	input N4END3;
	input NN4END0;
	input NN4END1;
	input NN4END2;
	input NN4END3;
	input bot2top0;
	input bot2top1;
	input bot2top2;
	input bot2top3;
	input bot2top4;
	input bot2top5;
	input bot2top6;
	input bot2top7;
	input bot2top8;
	input bot2top9;
	input E1END0;
	input E1END1;
	input E1END2;
	input E1END3;
	input E2MID0;
	input E2MID1;
	input E2MID2;
	input E2MID3;
	input E2MID4;
	input E2MID5;
	input E2MID6;
	input E2MID7;
	input E2END0;
	input E2END1;
	input E2END2;
	input E2END3;
	input E2END4;
	input E2END5;
	input E2END6;
	input E2END7;
	input EE4END0;
	input EE4END1;
	input EE4END2;
	input EE4END3;
	input E6END0;
	input E6END1;
	input S1END0;
	input S1END1;
	input S1END2;
	input S1END3;
	input S2MID0;
	input S2MID1;
	input S2MID2;
	input S2MID3;
	input S2MID4;
	input S2MID5;
	input S2MID6;
	input S2MID7;
	input S2END0;
	input S2END1;
	input S2END2;
	input S2END3;
	input S2END4;
	input S2END5;
	input S2END6;
	input S2END7;
	input S4END0;
	input S4END1;
	input S4END2;
	input S4END3;
	input SS4END0;
	input SS4END1;
	input SS4END2;
	input SS4END3;
	input W1END0;
	input W1END1;
	input W1END2;
	input W1END3;
	input W2MID0;
	input W2MID1;
	input W2MID2;
	input W2MID3;
	input W2MID4;
	input W2MID5;
	input W2MID6;
	input W2MID7;
	input W2END0;
	input W2END1;
	input W2END2;
	input W2END3;
	input W2END4;
	input W2END5;
	input W2END6;
	input W2END7;
	input WW4END0;
	input WW4END1;
	input WW4END2;
	input WW4END3;
	input W6END0;
	input W6END1;
	input J2MID_ABa_END0;
	input J2MID_ABa_END1;
	input J2MID_ABa_END2;
	input J2MID_ABa_END3;
	input J2MID_CDa_END0;
	input J2MID_CDa_END1;
	input J2MID_CDa_END2;
	input J2MID_CDa_END3;
	input J2MID_EFa_END0;
	input J2MID_EFa_END1;
	input J2MID_EFa_END2;
	input J2MID_EFa_END3;
	input J2MID_GHa_END0;
	input J2MID_GHa_END1;
	input J2MID_GHa_END2;
	input J2MID_GHa_END3;
	input J2MID_ABb_END0;
	input J2MID_ABb_END1;
	input J2MID_ABb_END2;
	input J2MID_ABb_END3;
	input J2MID_CDb_END0;
	input J2MID_CDb_END1;
	input J2MID_CDb_END2;
	input J2MID_CDb_END3;
	input J2MID_EFb_END0;
	input J2MID_EFb_END1;
	input J2MID_EFb_END2;
	input J2MID_EFb_END3;
	input J2MID_GHb_END0;
	input J2MID_GHb_END1;
	input J2MID_GHb_END2;
	input J2MID_GHb_END3;
	input J2END_AB_END0;
	input J2END_AB_END1;
	input J2END_AB_END2;
	input J2END_AB_END3;
	input J2END_CD_END0;
	input J2END_CD_END1;
	input J2END_CD_END2;
	input J2END_CD_END3;
	input J2END_EF_END0;
	input J2END_EF_END1;
	input J2END_EF_END2;
	input J2END_EF_END3;
	input J2END_GH_END0;
	input J2END_GH_END1;
	input J2END_GH_END2;
	input J2END_GH_END3;
	input JN2END0;
	input JN2END1;
	input JN2END2;
	input JN2END3;
	input JN2END4;
	input JN2END5;
	input JN2END6;
	input JN2END7;
	input JE2END0;
	input JE2END1;
	input JE2END2;
	input JE2END3;
	input JE2END4;
	input JE2END5;
	input JE2END6;
	input JE2END7;
	input JS2END0;
	input JS2END1;
	input JS2END2;
	input JS2END3;
	input JS2END4;
	input JS2END5;
	input JS2END6;
	input JS2END7;
	input JW2END0;
	input JW2END1;
	input JW2END2;
	input JW2END3;
	input JW2END4;
	input JW2END5;
	input JW2END6;
	input JW2END7;
	input J_l_AB_END0;
	input J_l_AB_END1;
	input J_l_AB_END2;
	input J_l_AB_END3;
	input J_l_CD_END0;
	input J_l_CD_END1;
	input J_l_CD_END2;
	input J_l_CD_END3;
	input J_l_EF_END0;
	input J_l_EF_END1;
	input J_l_EF_END2;
	input J_l_EF_END3;
	input J_l_GH_END0;
	input J_l_GH_END1;
	input J_l_GH_END2;
	input J_l_GH_END3;
	output N1BEG0;
	output N1BEG1;
	output N1BEG2;
	output N1BEG3;
	output N2BEG0;
	output N2BEG1;
	output N2BEG2;
	output N2BEG3;
	output N2BEG4;
	output N2BEG5;
	output N2BEG6;
	output N2BEG7;
	output N2BEGb0;
	output N2BEGb1;
	output N2BEGb2;
	output N2BEGb3;
	output N2BEGb4;
	output N2BEGb5;
	output N2BEGb6;
	output N2BEGb7;
	output N4BEG0;
	output N4BEG1;
	output N4BEG2;
	output N4BEG3;
	output NN4BEG0;
	output NN4BEG1;
	output NN4BEG2;
	output NN4BEG3;
	output E1BEG0;
	output E1BEG1;
	output E1BEG2;
	output E1BEG3;
	output E2BEG0;
	output E2BEG1;
	output E2BEG2;
	output E2BEG3;
	output E2BEG4;
	output E2BEG5;
	output E2BEG6;
	output E2BEG7;
	output E2BEGb0;
	output E2BEGb1;
	output E2BEGb2;
	output E2BEGb3;
	output E2BEGb4;
	output E2BEGb5;
	output E2BEGb6;
	output E2BEGb7;
	output EE4BEG0;
	output EE4BEG1;
	output EE4BEG2;
	output EE4BEG3;
	output E6BEG0;
	output E6BEG1;
	output S1BEG0;
	output S1BEG1;
	output S1BEG2;
	output S1BEG3;
	output S2BEG0;
	output S2BEG1;
	output S2BEG2;
	output S2BEG3;
	output S2BEG4;
	output S2BEG5;
	output S2BEG6;
	output S2BEG7;
	output S2BEGb0;
	output S2BEGb1;
	output S2BEGb2;
	output S2BEGb3;
	output S2BEGb4;
	output S2BEGb5;
	output S2BEGb6;
	output S2BEGb7;
	output S4BEG0;
	output S4BEG1;
	output S4BEG2;
	output S4BEG3;
	output SS4BEG0;
	output SS4BEG1;
	output SS4BEG2;
	output SS4BEG3;
	output top2bot0;
	output top2bot1;
	output top2bot2;
	output top2bot3;
	output top2bot4;
	output top2bot5;
	output top2bot6;
	output top2bot7;
	output top2bot8;
	output top2bot9;
	output top2bot10;
	output top2bot11;
	output top2bot12;
	output top2bot13;
	output top2bot14;
	output top2bot15;
	output top2bot16;
	output top2bot17;
	output W1BEG0;
	output W1BEG1;
	output W1BEG2;
	output W1BEG3;
	output W2BEG0;
	output W2BEG1;
	output W2BEG2;
	output W2BEG3;
	output W2BEG4;
	output W2BEG5;
	output W2BEG6;
	output W2BEG7;
	output W2BEGb0;
	output W2BEGb1;
	output W2BEGb2;
	output W2BEGb3;
	output W2BEGb4;
	output W2BEGb5;
	output W2BEGb6;
	output W2BEGb7;
	output WW4BEG0;
	output WW4BEG1;
	output WW4BEG2;
	output WW4BEG3;
	output W6BEG0;
	output W6BEG1;
	output J2MID_ABa_BEG0;
	output J2MID_ABa_BEG1;
	output J2MID_ABa_BEG2;
	output J2MID_ABa_BEG3;
	output J2MID_CDa_BEG0;
	output J2MID_CDa_BEG1;
	output J2MID_CDa_BEG2;
	output J2MID_CDa_BEG3;
	output J2MID_EFa_BEG0;
	output J2MID_EFa_BEG1;
	output J2MID_EFa_BEG2;
	output J2MID_EFa_BEG3;
	output J2MID_GHa_BEG0;
	output J2MID_GHa_BEG1;
	output J2MID_GHa_BEG2;
	output J2MID_GHa_BEG3;
	output J2MID_ABb_BEG0;
	output J2MID_ABb_BEG1;
	output J2MID_ABb_BEG2;
	output J2MID_ABb_BEG3;
	output J2MID_CDb_BEG0;
	output J2MID_CDb_BEG1;
	output J2MID_CDb_BEG2;
	output J2MID_CDb_BEG3;
	output J2MID_EFb_BEG0;
	output J2MID_EFb_BEG1;
	output J2MID_EFb_BEG2;
	output J2MID_EFb_BEG3;
	output J2MID_GHb_BEG0;
	output J2MID_GHb_BEG1;
	output J2MID_GHb_BEG2;
	output J2MID_GHb_BEG3;
	output J2END_AB_BEG0;
	output J2END_AB_BEG1;
	output J2END_AB_BEG2;
	output J2END_AB_BEG3;
	output J2END_CD_BEG0;
	output J2END_CD_BEG1;
	output J2END_CD_BEG2;
	output J2END_CD_BEG3;
	output J2END_EF_BEG0;
	output J2END_EF_BEG1;
	output J2END_EF_BEG2;
	output J2END_EF_BEG3;
	output J2END_GH_BEG0;
	output J2END_GH_BEG1;
	output J2END_GH_BEG2;
	output J2END_GH_BEG3;
	output JN2BEG0;
	output JN2BEG1;
	output JN2BEG2;
	output JN2BEG3;
	output JN2BEG4;
	output JN2BEG5;
	output JN2BEG6;
	output JN2BEG7;
	output JE2BEG0;
	output JE2BEG1;
	output JE2BEG2;
	output JE2BEG3;
	output JE2BEG4;
	output JE2BEG5;
	output JE2BEG6;
	output JE2BEG7;
	output JS2BEG0;
	output JS2BEG1;
	output JS2BEG2;
	output JS2BEG3;
	output JS2BEG4;
	output JS2BEG5;
	output JS2BEG6;
	output JS2BEG7;
	output JW2BEG0;
	output JW2BEG1;
	output JW2BEG2;
	output JW2BEG3;
	output JW2BEG4;
	output JW2BEG5;
	output JW2BEG6;
	output JW2BEG7;
	output J_l_AB_BEG0;
	output J_l_AB_BEG1;
	output J_l_AB_BEG2;
	output J_l_AB_BEG3;
	output J_l_CD_BEG0;
	output J_l_CD_BEG1;
	output J_l_CD_BEG2;
	output J_l_CD_BEG3;
	output J_l_EF_BEG0;
	output J_l_EF_BEG1;
	output J_l_EF_BEG2;
	output J_l_EF_BEG3;
	output J_l_GH_BEG0;
	output J_l_GH_BEG1;
	output J_l_GH_BEG2;
	output J_l_GH_BEG3;
	//global
	input [NoConfigBits-1:0] ConfigBits;
	input [NoConfigBits-1:0] ConfigBits_N;

	parameter GND0 = 1'b0;
	parameter GND = 1'b0;
	parameter VCC0 = 1'b1;
	parameter VCC = 1'b1;
	parameter VDD0 = 1'b1;
	parameter VDD = 1'b1;
	
	wire [4-1:0] N1BEG0_input;
	wire [4-1:0] N1BEG1_input;
	wire [4-1:0] N1BEG2_input;
	wire [4-1:0] N1BEG3_input;
	wire [1-1:0] N2BEG0_input;
	wire [1-1:0] N2BEG1_input;
	wire [1-1:0] N2BEG2_input;
	wire [1-1:0] N2BEG3_input;
	wire [1-1:0] N2BEG4_input;
	wire [1-1:0] N2BEG5_input;
	wire [1-1:0] N2BEG6_input;
	wire [1-1:0] N2BEG7_input;
	wire [1-1:0] N2BEGb0_input;
	wire [1-1:0] N2BEGb1_input;
	wire [1-1:0] N2BEGb2_input;
	wire [1-1:0] N2BEGb3_input;
	wire [1-1:0] N2BEGb4_input;
	wire [1-1:0] N2BEGb5_input;
	wire [1-1:0] N2BEGb6_input;
	wire [1-1:0] N2BEGb7_input;
	wire [4-1:0] N4BEG0_input;
	wire [4-1:0] N4BEG1_input;
	wire [4-1:0] N4BEG2_input;
	wire [4-1:0] N4BEG3_input;
	wire [8-1:0] NN4BEG0_input;
	wire [8-1:0] NN4BEG1_input;
	wire [8-1:0] NN4BEG2_input;
	wire [8-1:0] NN4BEG3_input;
	wire [4-1:0] E1BEG0_input;
	wire [4-1:0] E1BEG1_input;
	wire [4-1:0] E1BEG2_input;
	wire [4-1:0] E1BEG3_input;
	wire [1-1:0] E2BEG0_input;
	wire [1-1:0] E2BEG1_input;
	wire [1-1:0] E2BEG2_input;
	wire [1-1:0] E2BEG3_input;
	wire [1-1:0] E2BEG4_input;
	wire [1-1:0] E2BEG5_input;
	wire [1-1:0] E2BEG6_input;
	wire [1-1:0] E2BEG7_input;
	wire [1-1:0] E2BEGb0_input;
	wire [1-1:0] E2BEGb1_input;
	wire [1-1:0] E2BEGb2_input;
	wire [1-1:0] E2BEGb3_input;
	wire [1-1:0] E2BEGb4_input;
	wire [1-1:0] E2BEGb5_input;
	wire [1-1:0] E2BEGb6_input;
	wire [1-1:0] E2BEGb7_input;
	wire [8-1:0] EE4BEG0_input;
	wire [8-1:0] EE4BEG1_input;
	wire [8-1:0] EE4BEG2_input;
	wire [8-1:0] EE4BEG3_input;
	wire [16-1:0] E6BEG0_input;
	wire [16-1:0] E6BEG1_input;
	wire [4-1:0] S1BEG0_input;
	wire [4-1:0] S1BEG1_input;
	wire [4-1:0] S1BEG2_input;
	wire [4-1:0] S1BEG3_input;
	wire [1-1:0] S2BEG0_input;
	wire [1-1:0] S2BEG1_input;
	wire [1-1:0] S2BEG2_input;
	wire [1-1:0] S2BEG3_input;
	wire [1-1:0] S2BEG4_input;
	wire [1-1:0] S2BEG5_input;
	wire [1-1:0] S2BEG6_input;
	wire [1-1:0] S2BEG7_input;
	wire [1-1:0] S2BEGb0_input;
	wire [1-1:0] S2BEGb1_input;
	wire [1-1:0] S2BEGb2_input;
	wire [1-1:0] S2BEGb3_input;
	wire [1-1:0] S2BEGb4_input;
	wire [1-1:0] S2BEGb5_input;
	wire [1-1:0] S2BEGb6_input;
	wire [1-1:0] S2BEGb7_input;
	wire [4-1:0] S4BEG0_input;
	wire [4-1:0] S4BEG1_input;
	wire [4-1:0] S4BEG2_input;
	wire [4-1:0] S4BEG3_input;
	wire [8-1:0] SS4BEG0_input;
	wire [8-1:0] SS4BEG1_input;
	wire [8-1:0] SS4BEG2_input;
	wire [8-1:0] SS4BEG3_input;
	wire [4-1:0] top2bot0_input;
	wire [4-1:0] top2bot1_input;
	wire [4-1:0] top2bot2_input;
	wire [4-1:0] top2bot3_input;
	wire [4-1:0] top2bot4_input;
	wire [4-1:0] top2bot5_input;
	wire [4-1:0] top2bot6_input;
	wire [4-1:0] top2bot7_input;
	wire [4-1:0] top2bot8_input;
	wire [4-1:0] top2bot9_input;
	wire [4-1:0] top2bot10_input;
	wire [4-1:0] top2bot11_input;
	wire [4-1:0] top2bot12_input;
	wire [4-1:0] top2bot13_input;
	wire [4-1:0] top2bot14_input;
	wire [4-1:0] top2bot15_input;
	wire [8-1:0] top2bot16_input;
	wire [8-1:0] top2bot17_input;
	wire [4-1:0] W1BEG0_input;
	wire [4-1:0] W1BEG1_input;
	wire [4-1:0] W1BEG2_input;
	wire [4-1:0] W1BEG3_input;
	wire [1-1:0] W2BEG0_input;
	wire [1-1:0] W2BEG1_input;
	wire [1-1:0] W2BEG2_input;
	wire [1-1:0] W2BEG3_input;
	wire [1-1:0] W2BEG4_input;
	wire [1-1:0] W2BEG5_input;
	wire [1-1:0] W2BEG6_input;
	wire [1-1:0] W2BEG7_input;
	wire [1-1:0] W2BEGb0_input;
	wire [1-1:0] W2BEGb1_input;
	wire [1-1:0] W2BEGb2_input;
	wire [1-1:0] W2BEGb3_input;
	wire [1-1:0] W2BEGb4_input;
	wire [1-1:0] W2BEGb5_input;
	wire [1-1:0] W2BEGb6_input;
	wire [1-1:0] W2BEGb7_input;
	wire [8-1:0] WW4BEG0_input;
	wire [8-1:0] WW4BEG1_input;
	wire [8-1:0] WW4BEG2_input;
	wire [8-1:0] WW4BEG3_input;
	wire [16-1:0] W6BEG0_input;
	wire [16-1:0] W6BEG1_input;
	wire [4-1:0] J2MID_ABa_BEG0_input;
	wire [4-1:0] J2MID_ABa_BEG1_input;
	wire [4-1:0] J2MID_ABa_BEG2_input;
	wire [4-1:0] J2MID_ABa_BEG3_input;
	wire [4-1:0] J2MID_CDa_BEG0_input;
	wire [4-1:0] J2MID_CDa_BEG1_input;
	wire [4-1:0] J2MID_CDa_BEG2_input;
	wire [4-1:0] J2MID_CDa_BEG3_input;
	wire [4-1:0] J2MID_EFa_BEG0_input;
	wire [4-1:0] J2MID_EFa_BEG1_input;
	wire [4-1:0] J2MID_EFa_BEG2_input;
	wire [4-1:0] J2MID_EFa_BEG3_input;
	wire [4-1:0] J2MID_GHa_BEG0_input;
	wire [4-1:0] J2MID_GHa_BEG1_input;
	wire [4-1:0] J2MID_GHa_BEG2_input;
	wire [4-1:0] J2MID_GHa_BEG3_input;
	wire [4-1:0] J2MID_ABb_BEG0_input;
	wire [4-1:0] J2MID_ABb_BEG1_input;
	wire [4-1:0] J2MID_ABb_BEG2_input;
	wire [4-1:0] J2MID_ABb_BEG3_input;
	wire [4-1:0] J2MID_CDb_BEG0_input;
	wire [4-1:0] J2MID_CDb_BEG1_input;
	wire [4-1:0] J2MID_CDb_BEG2_input;
	wire [4-1:0] J2MID_CDb_BEG3_input;
	wire [4-1:0] J2MID_EFb_BEG0_input;
	wire [4-1:0] J2MID_EFb_BEG1_input;
	wire [4-1:0] J2MID_EFb_BEG2_input;
	wire [4-1:0] J2MID_EFb_BEG3_input;
	wire [4-1:0] J2MID_GHb_BEG0_input;
	wire [4-1:0] J2MID_GHb_BEG1_input;
	wire [4-1:0] J2MID_GHb_BEG2_input;
	wire [4-1:0] J2MID_GHb_BEG3_input;
	wire [4-1:0] J2END_AB_BEG0_input;
	wire [4-1:0] J2END_AB_BEG1_input;
	wire [4-1:0] J2END_AB_BEG2_input;
	wire [4-1:0] J2END_AB_BEG3_input;
	wire [4-1:0] J2END_CD_BEG0_input;
	wire [4-1:0] J2END_CD_BEG1_input;
	wire [4-1:0] J2END_CD_BEG2_input;
	wire [4-1:0] J2END_CD_BEG3_input;
	wire [4-1:0] J2END_EF_BEG0_input;
	wire [4-1:0] J2END_EF_BEG1_input;
	wire [4-1:0] J2END_EF_BEG2_input;
	wire [4-1:0] J2END_EF_BEG3_input;
	wire [4-1:0] J2END_GH_BEG0_input;
	wire [4-1:0] J2END_GH_BEG1_input;
	wire [4-1:0] J2END_GH_BEG2_input;
	wire [4-1:0] J2END_GH_BEG3_input;
	wire [16-1:0] JN2BEG0_input;
	wire [16-1:0] JN2BEG1_input;
	wire [16-1:0] JN2BEG2_input;
	wire [16-1:0] JN2BEG3_input;
	wire [16-1:0] JN2BEG4_input;
	wire [16-1:0] JN2BEG5_input;
	wire [16-1:0] JN2BEG6_input;
	wire [16-1:0] JN2BEG7_input;
	wire [16-1:0] JE2BEG0_input;
	wire [16-1:0] JE2BEG1_input;
	wire [16-1:0] JE2BEG2_input;
	wire [16-1:0] JE2BEG3_input;
	wire [16-1:0] JE2BEG4_input;
	wire [16-1:0] JE2BEG5_input;
	wire [16-1:0] JE2BEG6_input;
	wire [16-1:0] JE2BEG7_input;
	wire [16-1:0] JS2BEG0_input;
	wire [16-1:0] JS2BEG1_input;
	wire [16-1:0] JS2BEG2_input;
	wire [16-1:0] JS2BEG3_input;
	wire [16-1:0] JS2BEG4_input;
	wire [16-1:0] JS2BEG5_input;
	wire [16-1:0] JS2BEG6_input;
	wire [16-1:0] JS2BEG7_input;
	wire [16-1:0] JW2BEG0_input;
	wire [16-1:0] JW2BEG1_input;
	wire [16-1:0] JW2BEG2_input;
	wire [16-1:0] JW2BEG3_input;
	wire [16-1:0] JW2BEG4_input;
	wire [16-1:0] JW2BEG5_input;
	wire [16-1:0] JW2BEG6_input;
	wire [16-1:0] JW2BEG7_input;
	wire [4-1:0] J_l_AB_BEG0_input;
	wire [4-1:0] J_l_AB_BEG1_input;
	wire [4-1:0] J_l_AB_BEG2_input;
	wire [4-1:0] J_l_AB_BEG3_input;
	wire [4-1:0] J_l_CD_BEG0_input;
	wire [4-1:0] J_l_CD_BEG1_input;
	wire [4-1:0] J_l_CD_BEG2_input;
	wire [4-1:0] J_l_CD_BEG3_input;
	wire [4-1:0] J_l_EF_BEG0_input;
	wire [4-1:0] J_l_EF_BEG1_input;
	wire [4-1:0] J_l_EF_BEG2_input;
	wire [4-1:0] J_l_EF_BEG3_input;
	wire [4-1:0] J_l_GH_BEG0_input;
	wire [4-1:0] J_l_GH_BEG1_input;
	wire [4-1:0] J_l_GH_BEG2_input;
	wire [4-1:0] J_l_GH_BEG3_input;

	wire [2-1:0] DEBUG_select_N1BEG0;
	wire [2-1:0] DEBUG_select_N1BEG1;
	wire [2-1:0] DEBUG_select_N1BEG2;
	wire [2-1:0] DEBUG_select_N1BEG3;
	wire [2-1:0] DEBUG_select_N4BEG0;
	wire [2-1:0] DEBUG_select_N4BEG1;
	wire [2-1:0] DEBUG_select_N4BEG2;
	wire [2-1:0] DEBUG_select_N4BEG3;
	wire [3-1:0] DEBUG_select_NN4BEG0;
	wire [3-1:0] DEBUG_select_NN4BEG1;
	wire [3-1:0] DEBUG_select_NN4BEG2;
	wire [3-1:0] DEBUG_select_NN4BEG3;
	wire [2-1:0] DEBUG_select_E1BEG0;
	wire [2-1:0] DEBUG_select_E1BEG1;
	wire [2-1:0] DEBUG_select_E1BEG2;
	wire [2-1:0] DEBUG_select_E1BEG3;
	wire [3-1:0] DEBUG_select_EE4BEG0;
	wire [3-1:0] DEBUG_select_EE4BEG1;
	wire [3-1:0] DEBUG_select_EE4BEG2;
	wire [3-1:0] DEBUG_select_EE4BEG3;
	wire [4-1:0] DEBUG_select_E6BEG0;
	wire [4-1:0] DEBUG_select_E6BEG1;
	wire [2-1:0] DEBUG_select_S1BEG0;
	wire [2-1:0] DEBUG_select_S1BEG1;
	wire [2-1:0] DEBUG_select_S1BEG2;
	wire [2-1:0] DEBUG_select_S1BEG3;
	wire [2-1:0] DEBUG_select_S4BEG0;
	wire [2-1:0] DEBUG_select_S4BEG1;
	wire [2-1:0] DEBUG_select_S4BEG2;
	wire [2-1:0] DEBUG_select_S4BEG3;
	wire [3-1:0] DEBUG_select_SS4BEG0;
	wire [3-1:0] DEBUG_select_SS4BEG1;
	wire [3-1:0] DEBUG_select_SS4BEG2;
	wire [3-1:0] DEBUG_select_SS4BEG3;
	wire [2-1:0] DEBUG_select_top2bot0;
	wire [2-1:0] DEBUG_select_top2bot1;
	wire [2-1:0] DEBUG_select_top2bot2;
	wire [2-1:0] DEBUG_select_top2bot3;
	wire [2-1:0] DEBUG_select_top2bot4;
	wire [2-1:0] DEBUG_select_top2bot5;
	wire [2-1:0] DEBUG_select_top2bot6;
	wire [2-1:0] DEBUG_select_top2bot7;
	wire [2-1:0] DEBUG_select_top2bot8;
	wire [2-1:0] DEBUG_select_top2bot9;
	wire [2-1:0] DEBUG_select_top2bot10;
	wire [2-1:0] DEBUG_select_top2bot11;
	wire [2-1:0] DEBUG_select_top2bot12;
	wire [2-1:0] DEBUG_select_top2bot13;
	wire [2-1:0] DEBUG_select_top2bot14;
	wire [2-1:0] DEBUG_select_top2bot15;
	wire [3-1:0] DEBUG_select_top2bot16;
	wire [3-1:0] DEBUG_select_top2bot17;
	wire [2-1:0] DEBUG_select_W1BEG0;
	wire [2-1:0] DEBUG_select_W1BEG1;
	wire [2-1:0] DEBUG_select_W1BEG2;
	wire [2-1:0] DEBUG_select_W1BEG3;
	wire [3-1:0] DEBUG_select_WW4BEG0;
	wire [3-1:0] DEBUG_select_WW4BEG1;
	wire [3-1:0] DEBUG_select_WW4BEG2;
	wire [3-1:0] DEBUG_select_WW4BEG3;
	wire [4-1:0] DEBUG_select_W6BEG0;
	wire [4-1:0] DEBUG_select_W6BEG1;
	wire [2-1:0] DEBUG_select_J2MID_ABa_BEG0;
	wire [2-1:0] DEBUG_select_J2MID_ABa_BEG1;
	wire [2-1:0] DEBUG_select_J2MID_ABa_BEG2;
	wire [2-1:0] DEBUG_select_J2MID_ABa_BEG3;
	wire [2-1:0] DEBUG_select_J2MID_CDa_BEG0;
	wire [2-1:0] DEBUG_select_J2MID_CDa_BEG1;
	wire [2-1:0] DEBUG_select_J2MID_CDa_BEG2;
	wire [2-1:0] DEBUG_select_J2MID_CDa_BEG3;
	wire [2-1:0] DEBUG_select_J2MID_EFa_BEG0;
	wire [2-1:0] DEBUG_select_J2MID_EFa_BEG1;
	wire [2-1:0] DEBUG_select_J2MID_EFa_BEG2;
	wire [2-1:0] DEBUG_select_J2MID_EFa_BEG3;
	wire [2-1:0] DEBUG_select_J2MID_GHa_BEG0;
	wire [2-1:0] DEBUG_select_J2MID_GHa_BEG1;
	wire [2-1:0] DEBUG_select_J2MID_GHa_BEG2;
	wire [2-1:0] DEBUG_select_J2MID_GHa_BEG3;
	wire [2-1:0] DEBUG_select_J2MID_ABb_BEG0;
	wire [2-1:0] DEBUG_select_J2MID_ABb_BEG1;
	wire [2-1:0] DEBUG_select_J2MID_ABb_BEG2;
	wire [2-1:0] DEBUG_select_J2MID_ABb_BEG3;
	wire [2-1:0] DEBUG_select_J2MID_CDb_BEG0;
	wire [2-1:0] DEBUG_select_J2MID_CDb_BEG1;
	wire [2-1:0] DEBUG_select_J2MID_CDb_BEG2;
	wire [2-1:0] DEBUG_select_J2MID_CDb_BEG3;
	wire [2-1:0] DEBUG_select_J2MID_EFb_BEG0;
	wire [2-1:0] DEBUG_select_J2MID_EFb_BEG1;
	wire [2-1:0] DEBUG_select_J2MID_EFb_BEG2;
	wire [2-1:0] DEBUG_select_J2MID_EFb_BEG3;
	wire [2-1:0] DEBUG_select_J2MID_GHb_BEG0;
	wire [2-1:0] DEBUG_select_J2MID_GHb_BEG1;
	wire [2-1:0] DEBUG_select_J2MID_GHb_BEG2;
	wire [2-1:0] DEBUG_select_J2MID_GHb_BEG3;
	wire [2-1:0] DEBUG_select_J2END_AB_BEG0;
	wire [2-1:0] DEBUG_select_J2END_AB_BEG1;
	wire [2-1:0] DEBUG_select_J2END_AB_BEG2;
	wire [2-1:0] DEBUG_select_J2END_AB_BEG3;
	wire [2-1:0] DEBUG_select_J2END_CD_BEG0;
	wire [2-1:0] DEBUG_select_J2END_CD_BEG1;
	wire [2-1:0] DEBUG_select_J2END_CD_BEG2;
	wire [2-1:0] DEBUG_select_J2END_CD_BEG3;
	wire [2-1:0] DEBUG_select_J2END_EF_BEG0;
	wire [2-1:0] DEBUG_select_J2END_EF_BEG1;
	wire [2-1:0] DEBUG_select_J2END_EF_BEG2;
	wire [2-1:0] DEBUG_select_J2END_EF_BEG3;
	wire [2-1:0] DEBUG_select_J2END_GH_BEG0;
	wire [2-1:0] DEBUG_select_J2END_GH_BEG1;
	wire [2-1:0] DEBUG_select_J2END_GH_BEG2;
	wire [2-1:0] DEBUG_select_J2END_GH_BEG3;
	wire [4-1:0] DEBUG_select_JN2BEG0;
	wire [4-1:0] DEBUG_select_JN2BEG1;
	wire [4-1:0] DEBUG_select_JN2BEG2;
	wire [4-1:0] DEBUG_select_JN2BEG3;
	wire [4-1:0] DEBUG_select_JN2BEG4;
	wire [4-1:0] DEBUG_select_JN2BEG5;
	wire [4-1:0] DEBUG_select_JN2BEG6;
	wire [4-1:0] DEBUG_select_JN2BEG7;
	wire [4-1:0] DEBUG_select_JE2BEG0;
	wire [4-1:0] DEBUG_select_JE2BEG1;
	wire [4-1:0] DEBUG_select_JE2BEG2;
	wire [4-1:0] DEBUG_select_JE2BEG3;
	wire [4-1:0] DEBUG_select_JE2BEG4;
	wire [4-1:0] DEBUG_select_JE2BEG5;
	wire [4-1:0] DEBUG_select_JE2BEG6;
	wire [4-1:0] DEBUG_select_JE2BEG7;
	wire [4-1:0] DEBUG_select_JS2BEG0;
	wire [4-1:0] DEBUG_select_JS2BEG1;
	wire [4-1:0] DEBUG_select_JS2BEG2;
	wire [4-1:0] DEBUG_select_JS2BEG3;
	wire [4-1:0] DEBUG_select_JS2BEG4;
	wire [4-1:0] DEBUG_select_JS2BEG5;
	wire [4-1:0] DEBUG_select_JS2BEG6;
	wire [4-1:0] DEBUG_select_JS2BEG7;
	wire [4-1:0] DEBUG_select_JW2BEG0;
	wire [4-1:0] DEBUG_select_JW2BEG1;
	wire [4-1:0] DEBUG_select_JW2BEG2;
	wire [4-1:0] DEBUG_select_JW2BEG3;
	wire [4-1:0] DEBUG_select_JW2BEG4;
	wire [4-1:0] DEBUG_select_JW2BEG5;
	wire [4-1:0] DEBUG_select_JW2BEG6;
	wire [4-1:0] DEBUG_select_JW2BEG7;
	wire [2-1:0] DEBUG_select_J_l_AB_BEG0;
	wire [2-1:0] DEBUG_select_J_l_AB_BEG1;
	wire [2-1:0] DEBUG_select_J_l_AB_BEG2;
	wire [2-1:0] DEBUG_select_J_l_AB_BEG3;
	wire [2-1:0] DEBUG_select_J_l_CD_BEG0;
	wire [2-1:0] DEBUG_select_J_l_CD_BEG1;
	wire [2-1:0] DEBUG_select_J_l_CD_BEG2;
	wire [2-1:0] DEBUG_select_J_l_CD_BEG3;
	wire [2-1:0] DEBUG_select_J_l_EF_BEG0;
	wire [2-1:0] DEBUG_select_J_l_EF_BEG1;
	wire [2-1:0] DEBUG_select_J_l_EF_BEG2;
	wire [2-1:0] DEBUG_select_J_l_EF_BEG3;
	wire [2-1:0] DEBUG_select_J_l_GH_BEG0;
	wire [2-1:0] DEBUG_select_J_l_GH_BEG1;
	wire [2-1:0] DEBUG_select_J_l_GH_BEG2;
	wire [2-1:0] DEBUG_select_J_l_GH_BEG3;

// The configuration bits (if any) are just a long shift register

// This shift register is padded to an even number of flops/latches
// switch matrix multiplexer  N1BEG0 		MUX-4
	assign N1BEG0_input = {J_l_CD_END1,JW2END3,J2MID_CDb_END3,bot2top2};
	cus_mux41_buf inst_cus_mux41_buf_N1BEG0 (
	.A0 (N1BEG0_input[0]),
	.A1 (N1BEG0_input[1]),
	.A2 (N1BEG0_input[2]),
	.A3 (N1BEG0_input[3]),
	.S0 (ConfigBits[0+0]),
	.S0N (ConfigBits_N[0+0]),
	.S1 (ConfigBits[0+1]),
	.S1N (ConfigBits_N[0+1]),
	.X (N1BEG0)
	);

// switch matrix multiplexer  N1BEG1 		MUX-4
	assign N1BEG1_input = {J_l_EF_END2,JW2END0,J2MID_EFb_END0,bot2top3};
	cus_mux41_buf inst_cus_mux41_buf_N1BEG1 (
	.A0 (N1BEG1_input[0]),
	.A1 (N1BEG1_input[1]),
	.A2 (N1BEG1_input[2]),
	.A3 (N1BEG1_input[3]),
	.S0 (ConfigBits[2+0]),
	.S0N (ConfigBits_N[2+0]),
	.S1 (ConfigBits[2+1]),
	.S1N (ConfigBits_N[2+1]),
	.X (N1BEG1)
	);

// switch matrix multiplexer  N1BEG2 		MUX-4
	assign N1BEG2_input = {J_l_GH_END3,JW2END1,J2MID_GHb_END1,bot2top4};
	cus_mux41_buf inst_cus_mux41_buf_N1BEG2 (
	.A0 (N1BEG2_input[0]),
	.A1 (N1BEG2_input[1]),
	.A2 (N1BEG2_input[2]),
	.A3 (N1BEG2_input[3]),
	.S0 (ConfigBits[4+0]),
	.S0N (ConfigBits_N[4+0]),
	.S1 (ConfigBits[4+1]),
	.S1N (ConfigBits_N[4+1]),
	.X (N1BEG2)
	);

// switch matrix multiplexer  N1BEG3 		MUX-4
	assign N1BEG3_input = {J_l_AB_END0,JW2END2,J2MID_ABb_END2,bot2top5};
	cus_mux41_buf inst_cus_mux41_buf_N1BEG3 (
	.A0 (N1BEG3_input[0]),
	.A1 (N1BEG3_input[1]),
	.A2 (N1BEG3_input[2]),
	.A3 (N1BEG3_input[3]),
	.S0 (ConfigBits[6+0]),
	.S0N (ConfigBits_N[6+0]),
	.S1 (ConfigBits[6+1]),
	.S1N (ConfigBits_N[6+1]),
	.X (N1BEG3)
	);

// switch matrix multiplexer  N2BEG0 		MUX-1
	assign N2BEG0 = JN2END0;
// switch matrix multiplexer  N2BEG1 		MUX-1
	assign N2BEG1 = JN2END1;
// switch matrix multiplexer  N2BEG2 		MUX-1
	assign N2BEG2 = JN2END2;
// switch matrix multiplexer  N2BEG3 		MUX-1
	assign N2BEG3 = JN2END3;
// switch matrix multiplexer  N2BEG4 		MUX-1
	assign N2BEG4 = JN2END4;
// switch matrix multiplexer  N2BEG5 		MUX-1
	assign N2BEG5 = JN2END5;
// switch matrix multiplexer  N2BEG6 		MUX-1
	assign N2BEG6 = JN2END6;
// switch matrix multiplexer  N2BEG7 		MUX-1
	assign N2BEG7 = JN2END7;
// switch matrix multiplexer  N2BEGb0 		MUX-1
	assign N2BEGb0 = N2MID0;
// switch matrix multiplexer  N2BEGb1 		MUX-1
	assign N2BEGb1 = N2MID1;
// switch matrix multiplexer  N2BEGb2 		MUX-1
	assign N2BEGb2 = N2MID2;
// switch matrix multiplexer  N2BEGb3 		MUX-1
	assign N2BEGb3 = N2MID3;
// switch matrix multiplexer  N2BEGb4 		MUX-1
	assign N2BEGb4 = N2MID4;
// switch matrix multiplexer  N2BEGb5 		MUX-1
	assign N2BEGb5 = N2MID5;
// switch matrix multiplexer  N2BEGb6 		MUX-1
	assign N2BEGb6 = N2MID6;
// switch matrix multiplexer  N2BEGb7 		MUX-1
	assign N2BEGb7 = N2MID7;
// switch matrix multiplexer  N4BEG0 		MUX-4
	assign N4BEG0_input = {E6END1,bot2top4,N4END1,N2END2};
	cus_mux41_buf inst_cus_mux41_buf_N4BEG0 (
	.A0 (N4BEG0_input[0]),
	.A1 (N4BEG0_input[1]),
	.A2 (N4BEG0_input[2]),
	.A3 (N4BEG0_input[3]),
	.S0 (ConfigBits[8+0]),
	.S0N (ConfigBits_N[8+0]),
	.S1 (ConfigBits[8+1]),
	.S1N (ConfigBits_N[8+1]),
	.X (N4BEG0)
	);

// switch matrix multiplexer  N4BEG1 		MUX-4
	assign N4BEG1_input = {E6END0,bot2top5,N4END2,N2END3};
	cus_mux41_buf inst_cus_mux41_buf_N4BEG1 (
	.A0 (N4BEG1_input[0]),
	.A1 (N4BEG1_input[1]),
	.A2 (N4BEG1_input[2]),
	.A3 (N4BEG1_input[3]),
	.S0 (ConfigBits[10+0]),
	.S0N (ConfigBits_N[10+0]),
	.S1 (ConfigBits[10+1]),
	.S1N (ConfigBits_N[10+1]),
	.X (N4BEG1)
	);

// switch matrix multiplexer  N4BEG2 		MUX-4
	assign N4BEG2_input = {W6END1,bot2top6,N4END3,N2END0};
	cus_mux41_buf inst_cus_mux41_buf_N4BEG2 (
	.A0 (N4BEG2_input[0]),
	.A1 (N4BEG2_input[1]),
	.A2 (N4BEG2_input[2]),
	.A3 (N4BEG2_input[3]),
	.S0 (ConfigBits[12+0]),
	.S0N (ConfigBits_N[12+0]),
	.S1 (ConfigBits[12+1]),
	.S1N (ConfigBits_N[12+1]),
	.X (N4BEG2)
	);

// switch matrix multiplexer  N4BEG3 		MUX-4
	assign N4BEG3_input = {W6END0,bot2top7,N4END0,N2END1};
	cus_mux41_buf inst_cus_mux41_buf_N4BEG3 (
	.A0 (N4BEG3_input[0]),
	.A1 (N4BEG3_input[1]),
	.A2 (N4BEG3_input[2]),
	.A3 (N4BEG3_input[3]),
	.S0 (ConfigBits[14+0]),
	.S0N (ConfigBits_N[14+0]),
	.S1 (ConfigBits[14+1]),
	.S1N (ConfigBits_N[14+1]),
	.X (N4BEG3)
	);

// switch matrix multiplexer  NN4BEG0 		MUX-8
	assign NN4BEG0_input = {J2END_GH_END1,J2MID_CDb_END1,J2MID_ABb_END1,W1END2,E1END2,bot2top6,bot2top2,N1END2};
	cus_mux81_buf inst_cus_mux81_buf_NN4BEG0 (
	.A0 (NN4BEG0_input[0]),
	.A1 (NN4BEG0_input[1]),
	.A2 (NN4BEG0_input[2]),
	.A3 (NN4BEG0_input[3]),
	.A4 (NN4BEG0_input[4]),
	.A5 (NN4BEG0_input[5]),
	.A6 (NN4BEG0_input[6]),
	.A7 (NN4BEG0_input[7]),
	.S0 (ConfigBits[16+0]),
	.S0N (ConfigBits_N[16+0]),
	.S1 (ConfigBits[16+1]),
	.S1N (ConfigBits_N[16+1]),
	.S2 (ConfigBits[16+2]),
	.S2N (ConfigBits_N[16+2]),
	.X (NN4BEG0)
	);

// switch matrix multiplexer  NN4BEG1 		MUX-8
	assign NN4BEG1_input = {J2END_EF_END1,J2MID_CDa_END2,J2MID_ABa_END2,W1END3,E1END3,bot2top7,bot2top3,N1END3};
	cus_mux81_buf inst_cus_mux81_buf_NN4BEG1 (
	.A0 (NN4BEG1_input[0]),
	.A1 (NN4BEG1_input[1]),
	.A2 (NN4BEG1_input[2]),
	.A3 (NN4BEG1_input[3]),
	.A4 (NN4BEG1_input[4]),
	.A5 (NN4BEG1_input[5]),
	.A6 (NN4BEG1_input[6]),
	.A7 (NN4BEG1_input[7]),
	.S0 (ConfigBits[19+0]),
	.S0N (ConfigBits_N[19+0]),
	.S1 (ConfigBits[19+1]),
	.S1N (ConfigBits_N[19+1]),
	.S2 (ConfigBits[19+2]),
	.S2N (ConfigBits_N[19+2]),
	.X (NN4BEG1)
	);

// switch matrix multiplexer  NN4BEG2 		MUX-8
	assign NN4BEG2_input = {J2END_CD_END1,J2MID_GHb_END1,J2MID_EFb_END1,W1END0,E1END0,bot2top8,bot2top4,N1END0};
	cus_mux81_buf inst_cus_mux81_buf_NN4BEG2 (
	.A0 (NN4BEG2_input[0]),
	.A1 (NN4BEG2_input[1]),
	.A2 (NN4BEG2_input[2]),
	.A3 (NN4BEG2_input[3]),
	.A4 (NN4BEG2_input[4]),
	.A5 (NN4BEG2_input[5]),
	.A6 (NN4BEG2_input[6]),
	.A7 (NN4BEG2_input[7]),
	.S0 (ConfigBits[22+0]),
	.S0N (ConfigBits_N[22+0]),
	.S1 (ConfigBits[22+1]),
	.S1N (ConfigBits_N[22+1]),
	.S2 (ConfigBits[22+2]),
	.S2N (ConfigBits_N[22+2]),
	.X (NN4BEG2)
	);

// switch matrix multiplexer  NN4BEG3 		MUX-8
	assign NN4BEG3_input = {J2END_AB_END1,J2MID_GHa_END2,J2MID_EFa_END2,W1END1,E1END1,bot2top9,bot2top5,N1END1};
	cus_mux81_buf inst_cus_mux81_buf_NN4BEG3 (
	.A0 (NN4BEG3_input[0]),
	.A1 (NN4BEG3_input[1]),
	.A2 (NN4BEG3_input[2]),
	.A3 (NN4BEG3_input[3]),
	.A4 (NN4BEG3_input[4]),
	.A5 (NN4BEG3_input[5]),
	.A6 (NN4BEG3_input[6]),
	.A7 (NN4BEG3_input[7]),
	.S0 (ConfigBits[25+0]),
	.S0N (ConfigBits_N[25+0]),
	.S1 (ConfigBits[25+1]),
	.S1N (ConfigBits_N[25+1]),
	.S2 (ConfigBits[25+2]),
	.S2N (ConfigBits_N[25+2]),
	.X (NN4BEG3)
	);

// switch matrix multiplexer  E1BEG0 		MUX-4
	assign E1BEG0_input = {J_l_CD_END1,JN2END3,J2MID_CDb_END3,bot2top3};
	cus_mux41_buf inst_cus_mux41_buf_E1BEG0 (
	.A0 (E1BEG0_input[0]),
	.A1 (E1BEG0_input[1]),
	.A2 (E1BEG0_input[2]),
	.A3 (E1BEG0_input[3]),
	.S0 (ConfigBits[28+0]),
	.S0N (ConfigBits_N[28+0]),
	.S1 (ConfigBits[28+1]),
	.S1N (ConfigBits_N[28+1]),
	.X (E1BEG0)
	);

// switch matrix multiplexer  E1BEG1 		MUX-4
	assign E1BEG1_input = {J_l_EF_END2,JN2END0,J2MID_EFb_END0,bot2top4};
	cus_mux41_buf inst_cus_mux41_buf_E1BEG1 (
	.A0 (E1BEG1_input[0]),
	.A1 (E1BEG1_input[1]),
	.A2 (E1BEG1_input[2]),
	.A3 (E1BEG1_input[3]),
	.S0 (ConfigBits[30+0]),
	.S0N (ConfigBits_N[30+0]),
	.S1 (ConfigBits[30+1]),
	.S1N (ConfigBits_N[30+1]),
	.X (E1BEG1)
	);

// switch matrix multiplexer  E1BEG2 		MUX-4
	assign E1BEG2_input = {J_l_GH_END3,JN2END1,J2MID_GHb_END1,bot2top5};
	cus_mux41_buf inst_cus_mux41_buf_E1BEG2 (
	.A0 (E1BEG2_input[0]),
	.A1 (E1BEG2_input[1]),
	.A2 (E1BEG2_input[2]),
	.A3 (E1BEG2_input[3]),
	.S0 (ConfigBits[32+0]),
	.S0N (ConfigBits_N[32+0]),
	.S1 (ConfigBits[32+1]),
	.S1N (ConfigBits_N[32+1]),
	.X (E1BEG2)
	);

// switch matrix multiplexer  E1BEG3 		MUX-4
	assign E1BEG3_input = {J_l_AB_END0,JN2END2,J2MID_ABb_END2,bot2top6};
	cus_mux41_buf inst_cus_mux41_buf_E1BEG3 (
	.A0 (E1BEG3_input[0]),
	.A1 (E1BEG3_input[1]),
	.A2 (E1BEG3_input[2]),
	.A3 (E1BEG3_input[3]),
	.S0 (ConfigBits[34+0]),
	.S0N (ConfigBits_N[34+0]),
	.S1 (ConfigBits[34+1]),
	.S1N (ConfigBits_N[34+1]),
	.X (E1BEG3)
	);

// switch matrix multiplexer  E2BEG0 		MUX-1
	assign E2BEG0 = JE2END0;
// switch matrix multiplexer  E2BEG1 		MUX-1
	assign E2BEG1 = JE2END1;
// switch matrix multiplexer  E2BEG2 		MUX-1
	assign E2BEG2 = JE2END2;
// switch matrix multiplexer  E2BEG3 		MUX-1
	assign E2BEG3 = JE2END3;
// switch matrix multiplexer  E2BEG4 		MUX-1
	assign E2BEG4 = JE2END4;
// switch matrix multiplexer  E2BEG5 		MUX-1
	assign E2BEG5 = JE2END5;
// switch matrix multiplexer  E2BEG6 		MUX-1
	assign E2BEG6 = JE2END6;
// switch matrix multiplexer  E2BEG7 		MUX-1
	assign E2BEG7 = JE2END7;
// switch matrix multiplexer  E2BEGb0 		MUX-1
	assign E2BEGb0 = E2MID0;
// switch matrix multiplexer  E2BEGb1 		MUX-1
	assign E2BEGb1 = E2MID1;
// switch matrix multiplexer  E2BEGb2 		MUX-1
	assign E2BEGb2 = E2MID2;
// switch matrix multiplexer  E2BEGb3 		MUX-1
	assign E2BEGb3 = E2MID3;
// switch matrix multiplexer  E2BEGb4 		MUX-1
	assign E2BEGb4 = E2MID4;
// switch matrix multiplexer  E2BEGb5 		MUX-1
	assign E2BEGb5 = E2MID5;
// switch matrix multiplexer  E2BEGb6 		MUX-1
	assign E2BEGb6 = E2MID6;
// switch matrix multiplexer  E2BEGb7 		MUX-1
	assign E2BEGb7 = E2MID7;
// switch matrix multiplexer  EE4BEG0 		MUX-8
	assign EE4BEG0_input = {J2END_GH_END0,J2MID_CDb_END1,J2MID_ABb_END1,S1END2,E1END2,bot2top6,bot2top2,N1END2};
	cus_mux81_buf inst_cus_mux81_buf_EE4BEG0 (
	.A0 (EE4BEG0_input[0]),
	.A1 (EE4BEG0_input[1]),
	.A2 (EE4BEG0_input[2]),
	.A3 (EE4BEG0_input[3]),
	.A4 (EE4BEG0_input[4]),
	.A5 (EE4BEG0_input[5]),
	.A6 (EE4BEG0_input[6]),
	.A7 (EE4BEG0_input[7]),
	.S0 (ConfigBits[36+0]),
	.S0N (ConfigBits_N[36+0]),
	.S1 (ConfigBits[36+1]),
	.S1N (ConfigBits_N[36+1]),
	.S2 (ConfigBits[36+2]),
	.S2N (ConfigBits_N[36+2]),
	.X (EE4BEG0)
	);

// switch matrix multiplexer  EE4BEG1 		MUX-8
	assign EE4BEG1_input = {J2END_EF_END0,J2MID_CDa_END2,J2MID_ABa_END2,S1END3,E1END3,bot2top7,bot2top3,N1END3};
	cus_mux81_buf inst_cus_mux81_buf_EE4BEG1 (
	.A0 (EE4BEG1_input[0]),
	.A1 (EE4BEG1_input[1]),
	.A2 (EE4BEG1_input[2]),
	.A3 (EE4BEG1_input[3]),
	.A4 (EE4BEG1_input[4]),
	.A5 (EE4BEG1_input[5]),
	.A6 (EE4BEG1_input[6]),
	.A7 (EE4BEG1_input[7]),
	.S0 (ConfigBits[39+0]),
	.S0N (ConfigBits_N[39+0]),
	.S1 (ConfigBits[39+1]),
	.S1N (ConfigBits_N[39+1]),
	.S2 (ConfigBits[39+2]),
	.S2N (ConfigBits_N[39+2]),
	.X (EE4BEG1)
	);

// switch matrix multiplexer  EE4BEG2 		MUX-8
	assign EE4BEG2_input = {J2END_CD_END0,J2MID_GHb_END1,J2MID_EFb_END1,S1END0,E1END0,bot2top8,bot2top4,N1END0};
	cus_mux81_buf inst_cus_mux81_buf_EE4BEG2 (
	.A0 (EE4BEG2_input[0]),
	.A1 (EE4BEG2_input[1]),
	.A2 (EE4BEG2_input[2]),
	.A3 (EE4BEG2_input[3]),
	.A4 (EE4BEG2_input[4]),
	.A5 (EE4BEG2_input[5]),
	.A6 (EE4BEG2_input[6]),
	.A7 (EE4BEG2_input[7]),
	.S0 (ConfigBits[42+0]),
	.S0N (ConfigBits_N[42+0]),
	.S1 (ConfigBits[42+1]),
	.S1N (ConfigBits_N[42+1]),
	.S2 (ConfigBits[42+2]),
	.S2N (ConfigBits_N[42+2]),
	.X (EE4BEG2)
	);

// switch matrix multiplexer  EE4BEG3 		MUX-8
	assign EE4BEG3_input = {J2END_AB_END0,J2MID_GHa_END2,J2MID_EFa_END2,S1END1,E1END1,bot2top9,bot2top5,N1END1};
	cus_mux81_buf inst_cus_mux81_buf_EE4BEG3 (
	.A0 (EE4BEG3_input[0]),
	.A1 (EE4BEG3_input[1]),
	.A2 (EE4BEG3_input[2]),
	.A3 (EE4BEG3_input[3]),
	.A4 (EE4BEG3_input[4]),
	.A5 (EE4BEG3_input[5]),
	.A6 (EE4BEG3_input[6]),
	.A7 (EE4BEG3_input[7]),
	.S0 (ConfigBits[45+0]),
	.S0N (ConfigBits_N[45+0]),
	.S1 (ConfigBits[45+1]),
	.S1N (ConfigBits_N[45+1]),
	.S2 (ConfigBits[45+2]),
	.S2N (ConfigBits_N[45+2]),
	.X (EE4BEG3)
	);

// switch matrix multiplexer  E6BEG0 		MUX-16
	assign E6BEG0_input = {J2MID_GHb_END1,J2MID_EFb_END1,J2MID_CDb_END1,J2MID_ABb_END1,W1END3,E1END3,bot2top9,bot2top8,bot2top7,bot2top6,bot2top5,bot2top4,bot2top3,bot2top2,bot2top1,bot2top0};
	cus_mux161_buf inst_cus_mux161_buf_E6BEG0 (
	.A0 (E6BEG0_input[0]),
	.A1 (E6BEG0_input[1]),
	.A2 (E6BEG0_input[2]),
	.A3 (E6BEG0_input[3]),
	.A4 (E6BEG0_input[4]),
	.A5 (E6BEG0_input[5]),
	.A6 (E6BEG0_input[6]),
	.A7 (E6BEG0_input[7]),
	.A8 (E6BEG0_input[8]),
	.A9 (E6BEG0_input[9]),
	.A10 (E6BEG0_input[10]),
	.A11 (E6BEG0_input[11]),
	.A12 (E6BEG0_input[12]),
	.A13 (E6BEG0_input[13]),
	.A14 (E6BEG0_input[14]),
	.A15 (E6BEG0_input[15]),
	.S0 (ConfigBits[48+0]),
	.S0N (ConfigBits_N[48+0]),
	.S1 (ConfigBits[48+1]),
	.S1N (ConfigBits_N[48+1]),
	.S2 (ConfigBits[48+2]),
	.S2N (ConfigBits_N[48+2]),
	.S3 (ConfigBits[48+3]),
	.S3N (ConfigBits_N[48+3]),
	.X (E6BEG0)
	);

// switch matrix multiplexer  E6BEG1 		MUX-16
	assign E6BEG1_input = {J2MID_GHa_END2,J2MID_EFa_END2,J2MID_CDa_END2,J2MID_ABa_END2,W1END2,E1END2,bot2top9,bot2top8,bot2top7,bot2top6,bot2top5,bot2top4,bot2top3,bot2top2,bot2top1,bot2top0};
	cus_mux161_buf inst_cus_mux161_buf_E6BEG1 (
	.A0 (E6BEG1_input[0]),
	.A1 (E6BEG1_input[1]),
	.A2 (E6BEG1_input[2]),
	.A3 (E6BEG1_input[3]),
	.A4 (E6BEG1_input[4]),
	.A5 (E6BEG1_input[5]),
	.A6 (E6BEG1_input[6]),
	.A7 (E6BEG1_input[7]),
	.A8 (E6BEG1_input[8]),
	.A9 (E6BEG1_input[9]),
	.A10 (E6BEG1_input[10]),
	.A11 (E6BEG1_input[11]),
	.A12 (E6BEG1_input[12]),
	.A13 (E6BEG1_input[13]),
	.A14 (E6BEG1_input[14]),
	.A15 (E6BEG1_input[15]),
	.S0 (ConfigBits[52+0]),
	.S0N (ConfigBits_N[52+0]),
	.S1 (ConfigBits[52+1]),
	.S1N (ConfigBits_N[52+1]),
	.S2 (ConfigBits[52+2]),
	.S2N (ConfigBits_N[52+2]),
	.S3 (ConfigBits[52+3]),
	.S3N (ConfigBits_N[52+3]),
	.X (E6BEG1)
	);

// switch matrix multiplexer  S1BEG0 		MUX-4
	assign S1BEG0_input = {J_l_CD_END1,JE2END3,J2MID_CDb_END3,bot2top4};
	cus_mux41_buf inst_cus_mux41_buf_S1BEG0 (
	.A0 (S1BEG0_input[0]),
	.A1 (S1BEG0_input[1]),
	.A2 (S1BEG0_input[2]),
	.A3 (S1BEG0_input[3]),
	.S0 (ConfigBits[56+0]),
	.S0N (ConfigBits_N[56+0]),
	.S1 (ConfigBits[56+1]),
	.S1N (ConfigBits_N[56+1]),
	.X (S1BEG0)
	);

// switch matrix multiplexer  S1BEG1 		MUX-4
	assign S1BEG1_input = {J_l_EF_END2,JE2END0,J2MID_EFb_END0,bot2top5};
	cus_mux41_buf inst_cus_mux41_buf_S1BEG1 (
	.A0 (S1BEG1_input[0]),
	.A1 (S1BEG1_input[1]),
	.A2 (S1BEG1_input[2]),
	.A3 (S1BEG1_input[3]),
	.S0 (ConfigBits[58+0]),
	.S0N (ConfigBits_N[58+0]),
	.S1 (ConfigBits[58+1]),
	.S1N (ConfigBits_N[58+1]),
	.X (S1BEG1)
	);

// switch matrix multiplexer  S1BEG2 		MUX-4
	assign S1BEG2_input = {J_l_GH_END3,JE2END1,J2MID_GHb_END1,bot2top6};
	cus_mux41_buf inst_cus_mux41_buf_S1BEG2 (
	.A0 (S1BEG2_input[0]),
	.A1 (S1BEG2_input[1]),
	.A2 (S1BEG2_input[2]),
	.A3 (S1BEG2_input[3]),
	.S0 (ConfigBits[60+0]),
	.S0N (ConfigBits_N[60+0]),
	.S1 (ConfigBits[60+1]),
	.S1N (ConfigBits_N[60+1]),
	.X (S1BEG2)
	);

// switch matrix multiplexer  S1BEG3 		MUX-4
	assign S1BEG3_input = {J_l_AB_END0,JE2END2,J2MID_ABb_END2,bot2top7};
	cus_mux41_buf inst_cus_mux41_buf_S1BEG3 (
	.A0 (S1BEG3_input[0]),
	.A1 (S1BEG3_input[1]),
	.A2 (S1BEG3_input[2]),
	.A3 (S1BEG3_input[3]),
	.S0 (ConfigBits[62+0]),
	.S0N (ConfigBits_N[62+0]),
	.S1 (ConfigBits[62+1]),
	.S1N (ConfigBits_N[62+1]),
	.X (S1BEG3)
	);

// switch matrix multiplexer  S2BEG0 		MUX-1
	assign S2BEG0 = JS2END0;
// switch matrix multiplexer  S2BEG1 		MUX-1
	assign S2BEG1 = JS2END1;
// switch matrix multiplexer  S2BEG2 		MUX-1
	assign S2BEG2 = JS2END2;
// switch matrix multiplexer  S2BEG3 		MUX-1
	assign S2BEG3 = JS2END3;
// switch matrix multiplexer  S2BEG4 		MUX-1
	assign S2BEG4 = JS2END4;
// switch matrix multiplexer  S2BEG5 		MUX-1
	assign S2BEG5 = JS2END5;
// switch matrix multiplexer  S2BEG6 		MUX-1
	assign S2BEG6 = JS2END6;
// switch matrix multiplexer  S2BEG7 		MUX-1
	assign S2BEG7 = JS2END7;
// switch matrix multiplexer  S2BEGb0 		MUX-1
	assign S2BEGb0 = S2MID0;
// switch matrix multiplexer  S2BEGb1 		MUX-1
	assign S2BEGb1 = S2MID1;
// switch matrix multiplexer  S2BEGb2 		MUX-1
	assign S2BEGb2 = S2MID2;
// switch matrix multiplexer  S2BEGb3 		MUX-1
	assign S2BEGb3 = S2MID3;
// switch matrix multiplexer  S2BEGb4 		MUX-1
	assign S2BEGb4 = S2MID4;
// switch matrix multiplexer  S2BEGb5 		MUX-1
	assign S2BEGb5 = S2MID5;
// switch matrix multiplexer  S2BEGb6 		MUX-1
	assign S2BEGb6 = S2MID6;
// switch matrix multiplexer  S2BEGb7 		MUX-1
	assign S2BEGb7 = S2MID7;
// switch matrix multiplexer  S4BEG0 		MUX-4
	assign S4BEG0_input = {S4END1,S2END2,E6END1,bot2top0};
	cus_mux41_buf inst_cus_mux41_buf_S4BEG0 (
	.A0 (S4BEG0_input[0]),
	.A1 (S4BEG0_input[1]),
	.A2 (S4BEG0_input[2]),
	.A3 (S4BEG0_input[3]),
	.S0 (ConfigBits[64+0]),
	.S0N (ConfigBits_N[64+0]),
	.S1 (ConfigBits[64+1]),
	.S1N (ConfigBits_N[64+1]),
	.X (S4BEG0)
	);

// switch matrix multiplexer  S4BEG1 		MUX-4
	assign S4BEG1_input = {S4END2,S2END3,E6END0,bot2top1};
	cus_mux41_buf inst_cus_mux41_buf_S4BEG1 (
	.A0 (S4BEG1_input[0]),
	.A1 (S4BEG1_input[1]),
	.A2 (S4BEG1_input[2]),
	.A3 (S4BEG1_input[3]),
	.S0 (ConfigBits[66+0]),
	.S0N (ConfigBits_N[66+0]),
	.S1 (ConfigBits[66+1]),
	.S1N (ConfigBits_N[66+1]),
	.X (S4BEG1)
	);

// switch matrix multiplexer  S4BEG2 		MUX-4
	assign S4BEG2_input = {W6END1,S4END3,S2END0,bot2top2};
	cus_mux41_buf inst_cus_mux41_buf_S4BEG2 (
	.A0 (S4BEG2_input[0]),
	.A1 (S4BEG2_input[1]),
	.A2 (S4BEG2_input[2]),
	.A3 (S4BEG2_input[3]),
	.S0 (ConfigBits[68+0]),
	.S0N (ConfigBits_N[68+0]),
	.S1 (ConfigBits[68+1]),
	.S1N (ConfigBits_N[68+1]),
	.X (S4BEG2)
	);

// switch matrix multiplexer  S4BEG3 		MUX-4
	assign S4BEG3_input = {W6END0,S4END0,S2END1,bot2top3};
	cus_mux41_buf inst_cus_mux41_buf_S4BEG3 (
	.A0 (S4BEG3_input[0]),
	.A1 (S4BEG3_input[1]),
	.A2 (S4BEG3_input[2]),
	.A3 (S4BEG3_input[3]),
	.S0 (ConfigBits[70+0]),
	.S0N (ConfigBits_N[70+0]),
	.S1 (ConfigBits[70+1]),
	.S1N (ConfigBits_N[70+1]),
	.X (S4BEG3)
	);

// switch matrix multiplexer  SS4BEG0 		MUX-8
	assign SS4BEG0_input = {J2END_GH_END3,J2MID_CDb_END1,J2MID_ABb_END1,W1END2,E1END2,bot2top6,bot2top2,N1END2};
	cus_mux81_buf inst_cus_mux81_buf_SS4BEG0 (
	.A0 (SS4BEG0_input[0]),
	.A1 (SS4BEG0_input[1]),
	.A2 (SS4BEG0_input[2]),
	.A3 (SS4BEG0_input[3]),
	.A4 (SS4BEG0_input[4]),
	.A5 (SS4BEG0_input[5]),
	.A6 (SS4BEG0_input[6]),
	.A7 (SS4BEG0_input[7]),
	.S0 (ConfigBits[72+0]),
	.S0N (ConfigBits_N[72+0]),
	.S1 (ConfigBits[72+1]),
	.S1N (ConfigBits_N[72+1]),
	.S2 (ConfigBits[72+2]),
	.S2N (ConfigBits_N[72+2]),
	.X (SS4BEG0)
	);

// switch matrix multiplexer  SS4BEG1 		MUX-8
	assign SS4BEG1_input = {J2END_EF_END3,J2MID_CDa_END2,J2MID_ABa_END2,W1END3,E1END3,bot2top7,bot2top3,N1END3};
	cus_mux81_buf inst_cus_mux81_buf_SS4BEG1 (
	.A0 (SS4BEG1_input[0]),
	.A1 (SS4BEG1_input[1]),
	.A2 (SS4BEG1_input[2]),
	.A3 (SS4BEG1_input[3]),
	.A4 (SS4BEG1_input[4]),
	.A5 (SS4BEG1_input[5]),
	.A6 (SS4BEG1_input[6]),
	.A7 (SS4BEG1_input[7]),
	.S0 (ConfigBits[75+0]),
	.S0N (ConfigBits_N[75+0]),
	.S1 (ConfigBits[75+1]),
	.S1N (ConfigBits_N[75+1]),
	.S2 (ConfigBits[75+2]),
	.S2N (ConfigBits_N[75+2]),
	.X (SS4BEG1)
	);

// switch matrix multiplexer  SS4BEG2 		MUX-8
	assign SS4BEG2_input = {J2END_CD_END3,J2MID_GHb_END1,J2MID_EFb_END1,W1END0,E1END0,bot2top8,bot2top4,N1END0};
	cus_mux81_buf inst_cus_mux81_buf_SS4BEG2 (
	.A0 (SS4BEG2_input[0]),
	.A1 (SS4BEG2_input[1]),
	.A2 (SS4BEG2_input[2]),
	.A3 (SS4BEG2_input[3]),
	.A4 (SS4BEG2_input[4]),
	.A5 (SS4BEG2_input[5]),
	.A6 (SS4BEG2_input[6]),
	.A7 (SS4BEG2_input[7]),
	.S0 (ConfigBits[78+0]),
	.S0N (ConfigBits_N[78+0]),
	.S1 (ConfigBits[78+1]),
	.S1N (ConfigBits_N[78+1]),
	.S2 (ConfigBits[78+2]),
	.S2N (ConfigBits_N[78+2]),
	.X (SS4BEG2)
	);

// switch matrix multiplexer  SS4BEG3 		MUX-8
	assign SS4BEG3_input = {J2END_AB_END3,J2MID_GHa_END2,J2MID_EFa_END2,W1END1,E1END1,bot2top9,bot2top5,N1END1};
	cus_mux81_buf inst_cus_mux81_buf_SS4BEG3 (
	.A0 (SS4BEG3_input[0]),
	.A1 (SS4BEG3_input[1]),
	.A2 (SS4BEG3_input[2]),
	.A3 (SS4BEG3_input[3]),
	.A4 (SS4BEG3_input[4]),
	.A5 (SS4BEG3_input[5]),
	.A6 (SS4BEG3_input[6]),
	.A7 (SS4BEG3_input[7]),
	.S0 (ConfigBits[81+0]),
	.S0N (ConfigBits_N[81+0]),
	.S1 (ConfigBits[81+1]),
	.S1N (ConfigBits_N[81+1]),
	.S2 (ConfigBits[81+2]),
	.S2N (ConfigBits_N[81+2]),
	.X (SS4BEG3)
	);

// switch matrix multiplexer  top2bot0 		MUX-4
	assign top2bot0_input = {J_l_AB_END0,J2END_AB_END0,J2MID_ABb_END0,J2MID_ABa_END0};
	cus_mux41_buf inst_cus_mux41_buf_top2bot0 (
	.A0 (top2bot0_input[0]),
	.A1 (top2bot0_input[1]),
	.A2 (top2bot0_input[2]),
	.A3 (top2bot0_input[3]),
	.S0 (ConfigBits[84+0]),
	.S0N (ConfigBits_N[84+0]),
	.S1 (ConfigBits[84+1]),
	.S1N (ConfigBits_N[84+1]),
	.X (top2bot0)
	);

// switch matrix multiplexer  top2bot1 		MUX-4
	assign top2bot1_input = {J_l_AB_END1,J2END_AB_END1,J2MID_ABb_END1,J2MID_ABa_END1};
	cus_mux41_buf inst_cus_mux41_buf_top2bot1 (
	.A0 (top2bot1_input[0]),
	.A1 (top2bot1_input[1]),
	.A2 (top2bot1_input[2]),
	.A3 (top2bot1_input[3]),
	.S0 (ConfigBits[86+0]),
	.S0N (ConfigBits_N[86+0]),
	.S1 (ConfigBits[86+1]),
	.S1N (ConfigBits_N[86+1]),
	.X (top2bot1)
	);

// switch matrix multiplexer  top2bot2 		MUX-4
	assign top2bot2_input = {J_l_AB_END2,J2END_AB_END2,J2MID_ABb_END2,J2MID_ABa_END2};
	cus_mux41_buf inst_cus_mux41_buf_top2bot2 (
	.A0 (top2bot2_input[0]),
	.A1 (top2bot2_input[1]),
	.A2 (top2bot2_input[2]),
	.A3 (top2bot2_input[3]),
	.S0 (ConfigBits[88+0]),
	.S0N (ConfigBits_N[88+0]),
	.S1 (ConfigBits[88+1]),
	.S1N (ConfigBits_N[88+1]),
	.X (top2bot2)
	);

// switch matrix multiplexer  top2bot3 		MUX-4
	assign top2bot3_input = {J_l_AB_END3,J2END_AB_END3,J2MID_ABb_END3,J2MID_ABa_END3};
	cus_mux41_buf inst_cus_mux41_buf_top2bot3 (
	.A0 (top2bot3_input[0]),
	.A1 (top2bot3_input[1]),
	.A2 (top2bot3_input[2]),
	.A3 (top2bot3_input[3]),
	.S0 (ConfigBits[90+0]),
	.S0N (ConfigBits_N[90+0]),
	.S1 (ConfigBits[90+1]),
	.S1N (ConfigBits_N[90+1]),
	.X (top2bot3)
	);

// switch matrix multiplexer  top2bot4 		MUX-4
	assign top2bot4_input = {J_l_CD_END0,J2END_CD_END0,J2MID_CDb_END0,J2MID_CDa_END0};
	cus_mux41_buf inst_cus_mux41_buf_top2bot4 (
	.A0 (top2bot4_input[0]),
	.A1 (top2bot4_input[1]),
	.A2 (top2bot4_input[2]),
	.A3 (top2bot4_input[3]),
	.S0 (ConfigBits[92+0]),
	.S0N (ConfigBits_N[92+0]),
	.S1 (ConfigBits[92+1]),
	.S1N (ConfigBits_N[92+1]),
	.X (top2bot4)
	);

// switch matrix multiplexer  top2bot5 		MUX-4
	assign top2bot5_input = {J_l_CD_END1,J2END_CD_END1,J2MID_CDb_END1,J2MID_CDa_END1};
	cus_mux41_buf inst_cus_mux41_buf_top2bot5 (
	.A0 (top2bot5_input[0]),
	.A1 (top2bot5_input[1]),
	.A2 (top2bot5_input[2]),
	.A3 (top2bot5_input[3]),
	.S0 (ConfigBits[94+0]),
	.S0N (ConfigBits_N[94+0]),
	.S1 (ConfigBits[94+1]),
	.S1N (ConfigBits_N[94+1]),
	.X (top2bot5)
	);

// switch matrix multiplexer  top2bot6 		MUX-4
	assign top2bot6_input = {J_l_CD_END2,J2END_CD_END2,J2MID_CDb_END2,J2MID_CDa_END2};
	cus_mux41_buf inst_cus_mux41_buf_top2bot6 (
	.A0 (top2bot6_input[0]),
	.A1 (top2bot6_input[1]),
	.A2 (top2bot6_input[2]),
	.A3 (top2bot6_input[3]),
	.S0 (ConfigBits[96+0]),
	.S0N (ConfigBits_N[96+0]),
	.S1 (ConfigBits[96+1]),
	.S1N (ConfigBits_N[96+1]),
	.X (top2bot6)
	);

// switch matrix multiplexer  top2bot7 		MUX-4
	assign top2bot7_input = {J_l_CD_END3,J2END_CD_END3,J2MID_CDb_END3,J2MID_CDa_END3};
	cus_mux41_buf inst_cus_mux41_buf_top2bot7 (
	.A0 (top2bot7_input[0]),
	.A1 (top2bot7_input[1]),
	.A2 (top2bot7_input[2]),
	.A3 (top2bot7_input[3]),
	.S0 (ConfigBits[98+0]),
	.S0N (ConfigBits_N[98+0]),
	.S1 (ConfigBits[98+1]),
	.S1N (ConfigBits_N[98+1]),
	.X (top2bot7)
	);

// switch matrix multiplexer  top2bot8 		MUX-4
	assign top2bot8_input = {J_l_EF_END0,J2END_EF_END0,J2MID_EFb_END0,J2MID_EFa_END0};
	cus_mux41_buf inst_cus_mux41_buf_top2bot8 (
	.A0 (top2bot8_input[0]),
	.A1 (top2bot8_input[1]),
	.A2 (top2bot8_input[2]),
	.A3 (top2bot8_input[3]),
	.S0 (ConfigBits[100+0]),
	.S0N (ConfigBits_N[100+0]),
	.S1 (ConfigBits[100+1]),
	.S1N (ConfigBits_N[100+1]),
	.X (top2bot8)
	);

// switch matrix multiplexer  top2bot9 		MUX-4
	assign top2bot9_input = {J_l_EF_END1,J2END_EF_END1,J2MID_EFb_END1,J2MID_EFa_END1};
	cus_mux41_buf inst_cus_mux41_buf_top2bot9 (
	.A0 (top2bot9_input[0]),
	.A1 (top2bot9_input[1]),
	.A2 (top2bot9_input[2]),
	.A3 (top2bot9_input[3]),
	.S0 (ConfigBits[102+0]),
	.S0N (ConfigBits_N[102+0]),
	.S1 (ConfigBits[102+1]),
	.S1N (ConfigBits_N[102+1]),
	.X (top2bot9)
	);

// switch matrix multiplexer  top2bot10 		MUX-4
	assign top2bot10_input = {J_l_EF_END2,J2END_EF_END2,J2MID_EFb_END2,J2MID_EFa_END2};
	cus_mux41_buf inst_cus_mux41_buf_top2bot10 (
	.A0 (top2bot10_input[0]),
	.A1 (top2bot10_input[1]),
	.A2 (top2bot10_input[2]),
	.A3 (top2bot10_input[3]),
	.S0 (ConfigBits[104+0]),
	.S0N (ConfigBits_N[104+0]),
	.S1 (ConfigBits[104+1]),
	.S1N (ConfigBits_N[104+1]),
	.X (top2bot10)
	);

// switch matrix multiplexer  top2bot11 		MUX-4
	assign top2bot11_input = {J_l_EF_END3,J2END_EF_END3,J2MID_EFb_END3,J2MID_EFa_END3};
	cus_mux41_buf inst_cus_mux41_buf_top2bot11 (
	.A0 (top2bot11_input[0]),
	.A1 (top2bot11_input[1]),
	.A2 (top2bot11_input[2]),
	.A3 (top2bot11_input[3]),
	.S0 (ConfigBits[106+0]),
	.S0N (ConfigBits_N[106+0]),
	.S1 (ConfigBits[106+1]),
	.S1N (ConfigBits_N[106+1]),
	.X (top2bot11)
	);

// switch matrix multiplexer  top2bot12 		MUX-4
	assign top2bot12_input = {J_l_GH_END0,J2END_GH_END0,J2MID_GHb_END0,J2MID_GHa_END0};
	cus_mux41_buf inst_cus_mux41_buf_top2bot12 (
	.A0 (top2bot12_input[0]),
	.A1 (top2bot12_input[1]),
	.A2 (top2bot12_input[2]),
	.A3 (top2bot12_input[3]),
	.S0 (ConfigBits[108+0]),
	.S0N (ConfigBits_N[108+0]),
	.S1 (ConfigBits[108+1]),
	.S1N (ConfigBits_N[108+1]),
	.X (top2bot12)
	);

// switch matrix multiplexer  top2bot13 		MUX-4
	assign top2bot13_input = {J_l_GH_END1,J2END_GH_END1,J2MID_GHb_END1,J2MID_GHa_END1};
	cus_mux41_buf inst_cus_mux41_buf_top2bot13 (
	.A0 (top2bot13_input[0]),
	.A1 (top2bot13_input[1]),
	.A2 (top2bot13_input[2]),
	.A3 (top2bot13_input[3]),
	.S0 (ConfigBits[110+0]),
	.S0N (ConfigBits_N[110+0]),
	.S1 (ConfigBits[110+1]),
	.S1N (ConfigBits_N[110+1]),
	.X (top2bot13)
	);

// switch matrix multiplexer  top2bot14 		MUX-4
	assign top2bot14_input = {J_l_GH_END2,J2END_GH_END2,J2MID_GHb_END2,J2MID_GHa_END2};
	cus_mux41_buf inst_cus_mux41_buf_top2bot14 (
	.A0 (top2bot14_input[0]),
	.A1 (top2bot14_input[1]),
	.A2 (top2bot14_input[2]),
	.A3 (top2bot14_input[3]),
	.S0 (ConfigBits[112+0]),
	.S0N (ConfigBits_N[112+0]),
	.S1 (ConfigBits[112+1]),
	.S1N (ConfigBits_N[112+1]),
	.X (top2bot14)
	);

// switch matrix multiplexer  top2bot15 		MUX-4
	assign top2bot15_input = {J_l_GH_END3,J2END_GH_END3,J2MID_GHb_END3,J2MID_GHa_END3};
	cus_mux41_buf inst_cus_mux41_buf_top2bot15 (
	.A0 (top2bot15_input[0]),
	.A1 (top2bot15_input[1]),
	.A2 (top2bot15_input[2]),
	.A3 (top2bot15_input[3]),
	.S0 (ConfigBits[114+0]),
	.S0N (ConfigBits_N[114+0]),
	.S1 (ConfigBits[114+1]),
	.S1N (ConfigBits_N[114+1]),
	.X (top2bot15)
	);

// switch matrix multiplexer  top2bot16 		MUX-8
	assign top2bot16_input = {JW2END6,JW2END4,JS2END6,JS2END4,JE2END6,JE2END4,JN2END6,JN2END4};
	cus_mux81_buf inst_cus_mux81_buf_top2bot16 (
	.A0 (top2bot16_input[0]),
	.A1 (top2bot16_input[1]),
	.A2 (top2bot16_input[2]),
	.A3 (top2bot16_input[3]),
	.A4 (top2bot16_input[4]),
	.A5 (top2bot16_input[5]),
	.A6 (top2bot16_input[6]),
	.A7 (top2bot16_input[7]),
	.S0 (ConfigBits[116+0]),
	.S0N (ConfigBits_N[116+0]),
	.S1 (ConfigBits[116+1]),
	.S1N (ConfigBits_N[116+1]),
	.S2 (ConfigBits[116+2]),
	.S2N (ConfigBits_N[116+2]),
	.X (top2bot16)
	);

// switch matrix multiplexer  top2bot17 		MUX-8
	assign top2bot17_input = {JW2END7,JW2END5,JS2END7,JS2END5,JE2END7,JE2END5,JN2END7,JN2END5};
	cus_mux81_buf inst_cus_mux81_buf_top2bot17 (
	.A0 (top2bot17_input[0]),
	.A1 (top2bot17_input[1]),
	.A2 (top2bot17_input[2]),
	.A3 (top2bot17_input[3]),
	.A4 (top2bot17_input[4]),
	.A5 (top2bot17_input[5]),
	.A6 (top2bot17_input[6]),
	.A7 (top2bot17_input[7]),
	.S0 (ConfigBits[119+0]),
	.S0N (ConfigBits_N[119+0]),
	.S1 (ConfigBits[119+1]),
	.S1N (ConfigBits_N[119+1]),
	.S2 (ConfigBits[119+2]),
	.S2N (ConfigBits_N[119+2]),
	.X (top2bot17)
	);

// switch matrix multiplexer  W1BEG0 		MUX-4
	assign W1BEG0_input = {J_l_CD_END1,JS2END3,J2MID_CDb_END3,bot2top5};
	cus_mux41_buf inst_cus_mux41_buf_W1BEG0 (
	.A0 (W1BEG0_input[0]),
	.A1 (W1BEG0_input[1]),
	.A2 (W1BEG0_input[2]),
	.A3 (W1BEG0_input[3]),
	.S0 (ConfigBits[122+0]),
	.S0N (ConfigBits_N[122+0]),
	.S1 (ConfigBits[122+1]),
	.S1N (ConfigBits_N[122+1]),
	.X (W1BEG0)
	);

// switch matrix multiplexer  W1BEG1 		MUX-4
	assign W1BEG1_input = {J_l_EF_END2,JS2END0,J2MID_EFb_END0,bot2top6};
	cus_mux41_buf inst_cus_mux41_buf_W1BEG1 (
	.A0 (W1BEG1_input[0]),
	.A1 (W1BEG1_input[1]),
	.A2 (W1BEG1_input[2]),
	.A3 (W1BEG1_input[3]),
	.S0 (ConfigBits[124+0]),
	.S0N (ConfigBits_N[124+0]),
	.S1 (ConfigBits[124+1]),
	.S1N (ConfigBits_N[124+1]),
	.X (W1BEG1)
	);

// switch matrix multiplexer  W1BEG2 		MUX-4
	assign W1BEG2_input = {J_l_GH_END3,JS2END1,J2MID_GHb_END1,bot2top7};
	cus_mux41_buf inst_cus_mux41_buf_W1BEG2 (
	.A0 (W1BEG2_input[0]),
	.A1 (W1BEG2_input[1]),
	.A2 (W1BEG2_input[2]),
	.A3 (W1BEG2_input[3]),
	.S0 (ConfigBits[126+0]),
	.S0N (ConfigBits_N[126+0]),
	.S1 (ConfigBits[126+1]),
	.S1N (ConfigBits_N[126+1]),
	.X (W1BEG2)
	);

// switch matrix multiplexer  W1BEG3 		MUX-4
	assign W1BEG3_input = {J_l_AB_END0,JS2END2,J2MID_ABb_END2,bot2top0};
	cus_mux41_buf inst_cus_mux41_buf_W1BEG3 (
	.A0 (W1BEG3_input[0]),
	.A1 (W1BEG3_input[1]),
	.A2 (W1BEG3_input[2]),
	.A3 (W1BEG3_input[3]),
	.S0 (ConfigBits[128+0]),
	.S0N (ConfigBits_N[128+0]),
	.S1 (ConfigBits[128+1]),
	.S1N (ConfigBits_N[128+1]),
	.X (W1BEG3)
	);

// switch matrix multiplexer  W2BEG0 		MUX-1
	assign W2BEG0 = W2END0;
// switch matrix multiplexer  W2BEG1 		MUX-1
	assign W2BEG1 = JW2END1;
// switch matrix multiplexer  W2BEG2 		MUX-1
	assign W2BEG2 = JW2END2;
// switch matrix multiplexer  W2BEG3 		MUX-1
	assign W2BEG3 = W2END3;
// switch matrix multiplexer  W2BEG4 		MUX-1
	assign W2BEG4 = W2END4;
// switch matrix multiplexer  W2BEG5 		MUX-1
	assign W2BEG5 = JW2END5;
// switch matrix multiplexer  W2BEG6 		MUX-1
	assign W2BEG6 = JW2END6;
// switch matrix multiplexer  W2BEG7 		MUX-1
	assign W2BEG7 = W2END7;
// switch matrix multiplexer  W2BEGb0 		MUX-1
	assign W2BEGb0 = W2MID0;
// switch matrix multiplexer  W2BEGb1 		MUX-1
	assign W2BEGb1 = W2MID1;
// switch matrix multiplexer  W2BEGb2 		MUX-1
	assign W2BEGb2 = W2MID2;
// switch matrix multiplexer  W2BEGb3 		MUX-1
	assign W2BEGb3 = W2MID3;
// switch matrix multiplexer  W2BEGb4 		MUX-1
	assign W2BEGb4 = W2MID4;
// switch matrix multiplexer  W2BEGb5 		MUX-1
	assign W2BEGb5 = W2MID5;
// switch matrix multiplexer  W2BEGb6 		MUX-1
	assign W2BEGb6 = W2MID6;
// switch matrix multiplexer  W2BEGb7 		MUX-1
	assign W2BEGb7 = W2MID7;
// switch matrix multiplexer  WW4BEG0 		MUX-8
	assign WW4BEG0_input = {J2END_GH_END2,J2MID_CDb_END1,J2MID_ABb_END1,W1END2,S1END2,bot2top6,bot2top2,N1END2};
	cus_mux81_buf inst_cus_mux81_buf_WW4BEG0 (
	.A0 (WW4BEG0_input[0]),
	.A1 (WW4BEG0_input[1]),
	.A2 (WW4BEG0_input[2]),
	.A3 (WW4BEG0_input[3]),
	.A4 (WW4BEG0_input[4]),
	.A5 (WW4BEG0_input[5]),
	.A6 (WW4BEG0_input[6]),
	.A7 (WW4BEG0_input[7]),
	.S0 (ConfigBits[130+0]),
	.S0N (ConfigBits_N[130+0]),
	.S1 (ConfigBits[130+1]),
	.S1N (ConfigBits_N[130+1]),
	.S2 (ConfigBits[130+2]),
	.S2N (ConfigBits_N[130+2]),
	.X (WW4BEG0)
	);

// switch matrix multiplexer  WW4BEG1 		MUX-8
	assign WW4BEG1_input = {J2END_EF_END2,J2MID_CDa_END2,J2MID_ABa_END2,W1END3,S1END3,bot2top7,bot2top3,N1END3};
	cus_mux81_buf inst_cus_mux81_buf_WW4BEG1 (
	.A0 (WW4BEG1_input[0]),
	.A1 (WW4BEG1_input[1]),
	.A2 (WW4BEG1_input[2]),
	.A3 (WW4BEG1_input[3]),
	.A4 (WW4BEG1_input[4]),
	.A5 (WW4BEG1_input[5]),
	.A6 (WW4BEG1_input[6]),
	.A7 (WW4BEG1_input[7]),
	.S0 (ConfigBits[133+0]),
	.S0N (ConfigBits_N[133+0]),
	.S1 (ConfigBits[133+1]),
	.S1N (ConfigBits_N[133+1]),
	.S2 (ConfigBits[133+2]),
	.S2N (ConfigBits_N[133+2]),
	.X (WW4BEG1)
	);

// switch matrix multiplexer  WW4BEG2 		MUX-8
	assign WW4BEG2_input = {J2END_CD_END2,J2MID_GHb_END1,J2MID_EFb_END1,W1END0,S1END0,bot2top8,bot2top4,N1END0};
	cus_mux81_buf inst_cus_mux81_buf_WW4BEG2 (
	.A0 (WW4BEG2_input[0]),
	.A1 (WW4BEG2_input[1]),
	.A2 (WW4BEG2_input[2]),
	.A3 (WW4BEG2_input[3]),
	.A4 (WW4BEG2_input[4]),
	.A5 (WW4BEG2_input[5]),
	.A6 (WW4BEG2_input[6]),
	.A7 (WW4BEG2_input[7]),
	.S0 (ConfigBits[136+0]),
	.S0N (ConfigBits_N[136+0]),
	.S1 (ConfigBits[136+1]),
	.S1N (ConfigBits_N[136+1]),
	.S2 (ConfigBits[136+2]),
	.S2N (ConfigBits_N[136+2]),
	.X (WW4BEG2)
	);

// switch matrix multiplexer  WW4BEG3 		MUX-8
	assign WW4BEG3_input = {J2END_AB_END2,J2MID_GHa_END2,J2MID_EFa_END2,W1END1,S1END1,bot2top9,bot2top5,N1END1};
	cus_mux81_buf inst_cus_mux81_buf_WW4BEG3 (
	.A0 (WW4BEG3_input[0]),
	.A1 (WW4BEG3_input[1]),
	.A2 (WW4BEG3_input[2]),
	.A3 (WW4BEG3_input[3]),
	.A4 (WW4BEG3_input[4]),
	.A5 (WW4BEG3_input[5]),
	.A6 (WW4BEG3_input[6]),
	.A7 (WW4BEG3_input[7]),
	.S0 (ConfigBits[139+0]),
	.S0N (ConfigBits_N[139+0]),
	.S1 (ConfigBits[139+1]),
	.S1N (ConfigBits_N[139+1]),
	.S2 (ConfigBits[139+2]),
	.S2N (ConfigBits_N[139+2]),
	.X (WW4BEG3)
	);

// switch matrix multiplexer  W6BEG0 		MUX-16
	assign W6BEG0_input = {J2MID_GHb_END1,J2MID_EFb_END1,J2MID_CDb_END1,J2MID_ABb_END1,W1END3,E1END3,bot2top9,bot2top8,bot2top7,bot2top6,bot2top5,bot2top4,bot2top3,bot2top2,bot2top1,bot2top0};
	cus_mux161_buf inst_cus_mux161_buf_W6BEG0 (
	.A0 (W6BEG0_input[0]),
	.A1 (W6BEG0_input[1]),
	.A2 (W6BEG0_input[2]),
	.A3 (W6BEG0_input[3]),
	.A4 (W6BEG0_input[4]),
	.A5 (W6BEG0_input[5]),
	.A6 (W6BEG0_input[6]),
	.A7 (W6BEG0_input[7]),
	.A8 (W6BEG0_input[8]),
	.A9 (W6BEG0_input[9]),
	.A10 (W6BEG0_input[10]),
	.A11 (W6BEG0_input[11]),
	.A12 (W6BEG0_input[12]),
	.A13 (W6BEG0_input[13]),
	.A14 (W6BEG0_input[14]),
	.A15 (W6BEG0_input[15]),
	.S0 (ConfigBits[142+0]),
	.S0N (ConfigBits_N[142+0]),
	.S1 (ConfigBits[142+1]),
	.S1N (ConfigBits_N[142+1]),
	.S2 (ConfigBits[142+2]),
	.S2N (ConfigBits_N[142+2]),
	.S3 (ConfigBits[142+3]),
	.S3N (ConfigBits_N[142+3]),
	.X (W6BEG0)
	);

// switch matrix multiplexer  W6BEG1 		MUX-16
	assign W6BEG1_input = {J2MID_GHa_END2,J2MID_EFa_END2,J2MID_CDa_END2,J2MID_ABa_END2,W1END2,E1END2,bot2top9,bot2top8,bot2top7,bot2top6,bot2top5,bot2top4,bot2top3,bot2top2,bot2top1,bot2top0};
	cus_mux161_buf inst_cus_mux161_buf_W6BEG1 (
	.A0 (W6BEG1_input[0]),
	.A1 (W6BEG1_input[1]),
	.A2 (W6BEG1_input[2]),
	.A3 (W6BEG1_input[3]),
	.A4 (W6BEG1_input[4]),
	.A5 (W6BEG1_input[5]),
	.A6 (W6BEG1_input[6]),
	.A7 (W6BEG1_input[7]),
	.A8 (W6BEG1_input[8]),
	.A9 (W6BEG1_input[9]),
	.A10 (W6BEG1_input[10]),
	.A11 (W6BEG1_input[11]),
	.A12 (W6BEG1_input[12]),
	.A13 (W6BEG1_input[13]),
	.A14 (W6BEG1_input[14]),
	.A15 (W6BEG1_input[15]),
	.S0 (ConfigBits[146+0]),
	.S0N (ConfigBits_N[146+0]),
	.S1 (ConfigBits[146+1]),
	.S1N (ConfigBits_N[146+1]),
	.S2 (ConfigBits[146+2]),
	.S2N (ConfigBits_N[146+2]),
	.S3 (ConfigBits[146+3]),
	.S3N (ConfigBits_N[146+3]),
	.X (W6BEG1)
	);

// switch matrix multiplexer  J2MID_ABa_BEG0 		MUX-4
	assign J2MID_ABa_BEG0_input = {JN2END3,W2MID6,S2MID6,N2MID6};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_ABa_BEG0 (
	.A0 (J2MID_ABa_BEG0_input[0]),
	.A1 (J2MID_ABa_BEG0_input[1]),
	.A2 (J2MID_ABa_BEG0_input[2]),
	.A3 (J2MID_ABa_BEG0_input[3]),
	.S0 (ConfigBits[150+0]),
	.S0N (ConfigBits_N[150+0]),
	.S1 (ConfigBits[150+1]),
	.S1N (ConfigBits_N[150+1]),
	.X (J2MID_ABa_BEG0)
	);

// switch matrix multiplexer  J2MID_ABa_BEG1 		MUX-4
	assign J2MID_ABa_BEG1_input = {JE2END3,W2MID2,S2MID2,E2MID2};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_ABa_BEG1 (
	.A0 (J2MID_ABa_BEG1_input[0]),
	.A1 (J2MID_ABa_BEG1_input[1]),
	.A2 (J2MID_ABa_BEG1_input[2]),
	.A3 (J2MID_ABa_BEG1_input[3]),
	.S0 (ConfigBits[152+0]),
	.S0N (ConfigBits_N[152+0]),
	.S1 (ConfigBits[152+1]),
	.S1N (ConfigBits_N[152+1]),
	.X (J2MID_ABa_BEG1)
	);

// switch matrix multiplexer  J2MID_ABa_BEG2 		MUX-4
	assign J2MID_ABa_BEG2_input = {JS2END3,W2MID4,E2MID4,N2MID4};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_ABa_BEG2 (
	.A0 (J2MID_ABa_BEG2_input[0]),
	.A1 (J2MID_ABa_BEG2_input[1]),
	.A2 (J2MID_ABa_BEG2_input[2]),
	.A3 (J2MID_ABa_BEG2_input[3]),
	.S0 (ConfigBits[154+0]),
	.S0N (ConfigBits_N[154+0]),
	.S1 (ConfigBits[154+1]),
	.S1N (ConfigBits_N[154+1]),
	.X (J2MID_ABa_BEG2)
	);

// switch matrix multiplexer  J2MID_ABa_BEG3 		MUX-4
	assign J2MID_ABa_BEG3_input = {JW2END3,S2MID0,E2MID0,N2MID0};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_ABa_BEG3 (
	.A0 (J2MID_ABa_BEG3_input[0]),
	.A1 (J2MID_ABa_BEG3_input[1]),
	.A2 (J2MID_ABa_BEG3_input[2]),
	.A3 (J2MID_ABa_BEG3_input[3]),
	.S0 (ConfigBits[156+0]),
	.S0N (ConfigBits_N[156+0]),
	.S1 (ConfigBits[156+1]),
	.S1N (ConfigBits_N[156+1]),
	.X (J2MID_ABa_BEG3)
	);

// switch matrix multiplexer  J2MID_CDa_BEG0 		MUX-4
	assign J2MID_CDa_BEG0_input = {JN2END4,W2MID6,S2MID6,E2MID6};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_CDa_BEG0 (
	.A0 (J2MID_CDa_BEG0_input[0]),
	.A1 (J2MID_CDa_BEG0_input[1]),
	.A2 (J2MID_CDa_BEG0_input[2]),
	.A3 (J2MID_CDa_BEG0_input[3]),
	.S0 (ConfigBits[158+0]),
	.S0N (ConfigBits_N[158+0]),
	.S1 (ConfigBits[158+1]),
	.S1N (ConfigBits_N[158+1]),
	.X (J2MID_CDa_BEG0)
	);

// switch matrix multiplexer  J2MID_CDa_BEG1 		MUX-4
	assign J2MID_CDa_BEG1_input = {JE2END4,W2MID2,E2MID2,N2MID2};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_CDa_BEG1 (
	.A0 (J2MID_CDa_BEG1_input[0]),
	.A1 (J2MID_CDa_BEG1_input[1]),
	.A2 (J2MID_CDa_BEG1_input[2]),
	.A3 (J2MID_CDa_BEG1_input[3]),
	.S0 (ConfigBits[160+0]),
	.S0N (ConfigBits_N[160+0]),
	.S1 (ConfigBits[160+1]),
	.S1N (ConfigBits_N[160+1]),
	.X (J2MID_CDa_BEG1)
	);

// switch matrix multiplexer  J2MID_CDa_BEG2 		MUX-4
	assign J2MID_CDa_BEG2_input = {JS2END4,S2MID4,E2MID4,N2MID4};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_CDa_BEG2 (
	.A0 (J2MID_CDa_BEG2_input[0]),
	.A1 (J2MID_CDa_BEG2_input[1]),
	.A2 (J2MID_CDa_BEG2_input[2]),
	.A3 (J2MID_CDa_BEG2_input[3]),
	.S0 (ConfigBits[162+0]),
	.S0N (ConfigBits_N[162+0]),
	.S1 (ConfigBits[162+1]),
	.S1N (ConfigBits_N[162+1]),
	.X (J2MID_CDa_BEG2)
	);

// switch matrix multiplexer  J2MID_CDa_BEG3 		MUX-4
	assign J2MID_CDa_BEG3_input = {JW2END4,W2MID0,S2MID0,N2MID0};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_CDa_BEG3 (
	.A0 (J2MID_CDa_BEG3_input[0]),
	.A1 (J2MID_CDa_BEG3_input[1]),
	.A2 (J2MID_CDa_BEG3_input[2]),
	.A3 (J2MID_CDa_BEG3_input[3]),
	.S0 (ConfigBits[164+0]),
	.S0N (ConfigBits_N[164+0]),
	.S1 (ConfigBits[164+1]),
	.S1N (ConfigBits_N[164+1]),
	.X (J2MID_CDa_BEG3)
	);

// switch matrix multiplexer  J2MID_EFa_BEG0 		MUX-4
	assign J2MID_EFa_BEG0_input = {JN2END5,W2MID6,E2MID6,N2MID6};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_EFa_BEG0 (
	.A0 (J2MID_EFa_BEG0_input[0]),
	.A1 (J2MID_EFa_BEG0_input[1]),
	.A2 (J2MID_EFa_BEG0_input[2]),
	.A3 (J2MID_EFa_BEG0_input[3]),
	.S0 (ConfigBits[166+0]),
	.S0N (ConfigBits_N[166+0]),
	.S1 (ConfigBits[166+1]),
	.S1N (ConfigBits_N[166+1]),
	.X (J2MID_EFa_BEG0)
	);

// switch matrix multiplexer  J2MID_EFa_BEG1 		MUX-4
	assign J2MID_EFa_BEG1_input = {JE2END5,S2MID2,E2MID2,N2MID2};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_EFa_BEG1 (
	.A0 (J2MID_EFa_BEG1_input[0]),
	.A1 (J2MID_EFa_BEG1_input[1]),
	.A2 (J2MID_EFa_BEG1_input[2]),
	.A3 (J2MID_EFa_BEG1_input[3]),
	.S0 (ConfigBits[168+0]),
	.S0N (ConfigBits_N[168+0]),
	.S1 (ConfigBits[168+1]),
	.S1N (ConfigBits_N[168+1]),
	.X (J2MID_EFa_BEG1)
	);

// switch matrix multiplexer  J2MID_EFa_BEG2 		MUX-4
	assign J2MID_EFa_BEG2_input = {JS2END5,W2MID4,S2MID4,N2MID4};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_EFa_BEG2 (
	.A0 (J2MID_EFa_BEG2_input[0]),
	.A1 (J2MID_EFa_BEG2_input[1]),
	.A2 (J2MID_EFa_BEG2_input[2]),
	.A3 (J2MID_EFa_BEG2_input[3]),
	.S0 (ConfigBits[170+0]),
	.S0N (ConfigBits_N[170+0]),
	.S1 (ConfigBits[170+1]),
	.S1N (ConfigBits_N[170+1]),
	.X (J2MID_EFa_BEG2)
	);

// switch matrix multiplexer  J2MID_EFa_BEG3 		MUX-4
	assign J2MID_EFa_BEG3_input = {JW2END5,W2MID0,S2MID0,E2MID0};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_EFa_BEG3 (
	.A0 (J2MID_EFa_BEG3_input[0]),
	.A1 (J2MID_EFa_BEG3_input[1]),
	.A2 (J2MID_EFa_BEG3_input[2]),
	.A3 (J2MID_EFa_BEG3_input[3]),
	.S0 (ConfigBits[172+0]),
	.S0N (ConfigBits_N[172+0]),
	.S1 (ConfigBits[172+1]),
	.S1N (ConfigBits_N[172+1]),
	.X (J2MID_EFa_BEG3)
	);

// switch matrix multiplexer  J2MID_GHa_BEG0 		MUX-4
	assign J2MID_GHa_BEG0_input = {JN2END6,S2MID6,E2MID6,N2MID6};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_GHa_BEG0 (
	.A0 (J2MID_GHa_BEG0_input[0]),
	.A1 (J2MID_GHa_BEG0_input[1]),
	.A2 (J2MID_GHa_BEG0_input[2]),
	.A3 (J2MID_GHa_BEG0_input[3]),
	.S0 (ConfigBits[174+0]),
	.S0N (ConfigBits_N[174+0]),
	.S1 (ConfigBits[174+1]),
	.S1N (ConfigBits_N[174+1]),
	.X (J2MID_GHa_BEG0)
	);

// switch matrix multiplexer  J2MID_GHa_BEG1 		MUX-4
	assign J2MID_GHa_BEG1_input = {JE2END6,W2MID2,S2MID2,N2MID2};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_GHa_BEG1 (
	.A0 (J2MID_GHa_BEG1_input[0]),
	.A1 (J2MID_GHa_BEG1_input[1]),
	.A2 (J2MID_GHa_BEG1_input[2]),
	.A3 (J2MID_GHa_BEG1_input[3]),
	.S0 (ConfigBits[176+0]),
	.S0N (ConfigBits_N[176+0]),
	.S1 (ConfigBits[176+1]),
	.S1N (ConfigBits_N[176+1]),
	.X (J2MID_GHa_BEG1)
	);

// switch matrix multiplexer  J2MID_GHa_BEG2 		MUX-4
	assign J2MID_GHa_BEG2_input = {JS2END6,W2MID4,S2MID4,E2MID4};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_GHa_BEG2 (
	.A0 (J2MID_GHa_BEG2_input[0]),
	.A1 (J2MID_GHa_BEG2_input[1]),
	.A2 (J2MID_GHa_BEG2_input[2]),
	.A3 (J2MID_GHa_BEG2_input[3]),
	.S0 (ConfigBits[178+0]),
	.S0N (ConfigBits_N[178+0]),
	.S1 (ConfigBits[178+1]),
	.S1N (ConfigBits_N[178+1]),
	.X (J2MID_GHa_BEG2)
	);

// switch matrix multiplexer  J2MID_GHa_BEG3 		MUX-4
	assign J2MID_GHa_BEG3_input = {JW2END6,W2MID0,E2MID0,N2MID0};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_GHa_BEG3 (
	.A0 (J2MID_GHa_BEG3_input[0]),
	.A1 (J2MID_GHa_BEG3_input[1]),
	.A2 (J2MID_GHa_BEG3_input[2]),
	.A3 (J2MID_GHa_BEG3_input[3]),
	.S0 (ConfigBits[180+0]),
	.S0N (ConfigBits_N[180+0]),
	.S1 (ConfigBits[180+1]),
	.S1N (ConfigBits_N[180+1]),
	.X (J2MID_GHa_BEG3)
	);

// switch matrix multiplexer  J2MID_ABb_BEG0 		MUX-4
	assign J2MID_ABb_BEG0_input = {W2MID7,S2MID7,E2MID7,N2MID7};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_ABb_BEG0 (
	.A0 (J2MID_ABb_BEG0_input[0]),
	.A1 (J2MID_ABb_BEG0_input[1]),
	.A2 (J2MID_ABb_BEG0_input[2]),
	.A3 (J2MID_ABb_BEG0_input[3]),
	.S0 (ConfigBits[182+0]),
	.S0N (ConfigBits_N[182+0]),
	.S1 (ConfigBits[182+1]),
	.S1N (ConfigBits_N[182+1]),
	.X (J2MID_ABb_BEG0)
	);

// switch matrix multiplexer  J2MID_ABb_BEG1 		MUX-4
	assign J2MID_ABb_BEG1_input = {W2MID3,S2MID3,E2MID3,N2MID3};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_ABb_BEG1 (
	.A0 (J2MID_ABb_BEG1_input[0]),
	.A1 (J2MID_ABb_BEG1_input[1]),
	.A2 (J2MID_ABb_BEG1_input[2]),
	.A3 (J2MID_ABb_BEG1_input[3]),
	.S0 (ConfigBits[184+0]),
	.S0N (ConfigBits_N[184+0]),
	.S1 (ConfigBits[184+1]),
	.S1N (ConfigBits_N[184+1]),
	.X (J2MID_ABb_BEG1)
	);

// switch matrix multiplexer  J2MID_ABb_BEG2 		MUX-4
	assign J2MID_ABb_BEG2_input = {W2MID5,S2MID5,E2MID5,N2MID5};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_ABb_BEG2 (
	.A0 (J2MID_ABb_BEG2_input[0]),
	.A1 (J2MID_ABb_BEG2_input[1]),
	.A2 (J2MID_ABb_BEG2_input[2]),
	.A3 (J2MID_ABb_BEG2_input[3]),
	.S0 (ConfigBits[186+0]),
	.S0N (ConfigBits_N[186+0]),
	.S1 (ConfigBits[186+1]),
	.S1N (ConfigBits_N[186+1]),
	.X (J2MID_ABb_BEG2)
	);

// switch matrix multiplexer  J2MID_ABb_BEG3 		MUX-4
	assign J2MID_ABb_BEG3_input = {W2MID1,S2MID1,E2MID1,N2MID1};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_ABb_BEG3 (
	.A0 (J2MID_ABb_BEG3_input[0]),
	.A1 (J2MID_ABb_BEG3_input[1]),
	.A2 (J2MID_ABb_BEG3_input[2]),
	.A3 (J2MID_ABb_BEG3_input[3]),
	.S0 (ConfigBits[188+0]),
	.S0N (ConfigBits_N[188+0]),
	.S1 (ConfigBits[188+1]),
	.S1N (ConfigBits_N[188+1]),
	.X (J2MID_ABb_BEG3)
	);

// switch matrix multiplexer  J2MID_CDb_BEG0 		MUX-4
	assign J2MID_CDb_BEG0_input = {W2MID7,S2MID7,E2MID7,N2MID7};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_CDb_BEG0 (
	.A0 (J2MID_CDb_BEG0_input[0]),
	.A1 (J2MID_CDb_BEG0_input[1]),
	.A2 (J2MID_CDb_BEG0_input[2]),
	.A3 (J2MID_CDb_BEG0_input[3]),
	.S0 (ConfigBits[190+0]),
	.S0N (ConfigBits_N[190+0]),
	.S1 (ConfigBits[190+1]),
	.S1N (ConfigBits_N[190+1]),
	.X (J2MID_CDb_BEG0)
	);

// switch matrix multiplexer  J2MID_CDb_BEG1 		MUX-4
	assign J2MID_CDb_BEG1_input = {W2MID3,S2MID3,E2MID3,N2MID3};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_CDb_BEG1 (
	.A0 (J2MID_CDb_BEG1_input[0]),
	.A1 (J2MID_CDb_BEG1_input[1]),
	.A2 (J2MID_CDb_BEG1_input[2]),
	.A3 (J2MID_CDb_BEG1_input[3]),
	.S0 (ConfigBits[192+0]),
	.S0N (ConfigBits_N[192+0]),
	.S1 (ConfigBits[192+1]),
	.S1N (ConfigBits_N[192+1]),
	.X (J2MID_CDb_BEG1)
	);

// switch matrix multiplexer  J2MID_CDb_BEG2 		MUX-4
	assign J2MID_CDb_BEG2_input = {W2MID5,S2MID5,E2MID5,N2MID5};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_CDb_BEG2 (
	.A0 (J2MID_CDb_BEG2_input[0]),
	.A1 (J2MID_CDb_BEG2_input[1]),
	.A2 (J2MID_CDb_BEG2_input[2]),
	.A3 (J2MID_CDb_BEG2_input[3]),
	.S0 (ConfigBits[194+0]),
	.S0N (ConfigBits_N[194+0]),
	.S1 (ConfigBits[194+1]),
	.S1N (ConfigBits_N[194+1]),
	.X (J2MID_CDb_BEG2)
	);

// switch matrix multiplexer  J2MID_CDb_BEG3 		MUX-4
	assign J2MID_CDb_BEG3_input = {W2MID1,S2MID1,E2MID1,N2MID1};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_CDb_BEG3 (
	.A0 (J2MID_CDb_BEG3_input[0]),
	.A1 (J2MID_CDb_BEG3_input[1]),
	.A2 (J2MID_CDb_BEG3_input[2]),
	.A3 (J2MID_CDb_BEG3_input[3]),
	.S0 (ConfigBits[196+0]),
	.S0N (ConfigBits_N[196+0]),
	.S1 (ConfigBits[196+1]),
	.S1N (ConfigBits_N[196+1]),
	.X (J2MID_CDb_BEG3)
	);

// switch matrix multiplexer  J2MID_EFb_BEG0 		MUX-4
	assign J2MID_EFb_BEG0_input = {W2MID7,S2MID7,E2MID7,N2MID7};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_EFb_BEG0 (
	.A0 (J2MID_EFb_BEG0_input[0]),
	.A1 (J2MID_EFb_BEG0_input[1]),
	.A2 (J2MID_EFb_BEG0_input[2]),
	.A3 (J2MID_EFb_BEG0_input[3]),
	.S0 (ConfigBits[198+0]),
	.S0N (ConfigBits_N[198+0]),
	.S1 (ConfigBits[198+1]),
	.S1N (ConfigBits_N[198+1]),
	.X (J2MID_EFb_BEG0)
	);

// switch matrix multiplexer  J2MID_EFb_BEG1 		MUX-4
	assign J2MID_EFb_BEG1_input = {W2MID3,S2MID3,E2MID3,N2MID3};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_EFb_BEG1 (
	.A0 (J2MID_EFb_BEG1_input[0]),
	.A1 (J2MID_EFb_BEG1_input[1]),
	.A2 (J2MID_EFb_BEG1_input[2]),
	.A3 (J2MID_EFb_BEG1_input[3]),
	.S0 (ConfigBits[200+0]),
	.S0N (ConfigBits_N[200+0]),
	.S1 (ConfigBits[200+1]),
	.S1N (ConfigBits_N[200+1]),
	.X (J2MID_EFb_BEG1)
	);

// switch matrix multiplexer  J2MID_EFb_BEG2 		MUX-4
	assign J2MID_EFb_BEG2_input = {W2MID5,S2MID5,E2MID5,N2MID5};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_EFb_BEG2 (
	.A0 (J2MID_EFb_BEG2_input[0]),
	.A1 (J2MID_EFb_BEG2_input[1]),
	.A2 (J2MID_EFb_BEG2_input[2]),
	.A3 (J2MID_EFb_BEG2_input[3]),
	.S0 (ConfigBits[202+0]),
	.S0N (ConfigBits_N[202+0]),
	.S1 (ConfigBits[202+1]),
	.S1N (ConfigBits_N[202+1]),
	.X (J2MID_EFb_BEG2)
	);

// switch matrix multiplexer  J2MID_EFb_BEG3 		MUX-4
	assign J2MID_EFb_BEG3_input = {W2MID1,S2MID1,E2MID1,N2MID1};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_EFb_BEG3 (
	.A0 (J2MID_EFb_BEG3_input[0]),
	.A1 (J2MID_EFb_BEG3_input[1]),
	.A2 (J2MID_EFb_BEG3_input[2]),
	.A3 (J2MID_EFb_BEG3_input[3]),
	.S0 (ConfigBits[204+0]),
	.S0N (ConfigBits_N[204+0]),
	.S1 (ConfigBits[204+1]),
	.S1N (ConfigBits_N[204+1]),
	.X (J2MID_EFb_BEG3)
	);

// switch matrix multiplexer  J2MID_GHb_BEG0 		MUX-4
	assign J2MID_GHb_BEG0_input = {W2MID7,S2MID7,E2MID7,N2MID7};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_GHb_BEG0 (
	.A0 (J2MID_GHb_BEG0_input[0]),
	.A1 (J2MID_GHb_BEG0_input[1]),
	.A2 (J2MID_GHb_BEG0_input[2]),
	.A3 (J2MID_GHb_BEG0_input[3]),
	.S0 (ConfigBits[206+0]),
	.S0N (ConfigBits_N[206+0]),
	.S1 (ConfigBits[206+1]),
	.S1N (ConfigBits_N[206+1]),
	.X (J2MID_GHb_BEG0)
	);

// switch matrix multiplexer  J2MID_GHb_BEG1 		MUX-4
	assign J2MID_GHb_BEG1_input = {W2MID3,S2MID3,E2MID3,N2MID3};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_GHb_BEG1 (
	.A0 (J2MID_GHb_BEG1_input[0]),
	.A1 (J2MID_GHb_BEG1_input[1]),
	.A2 (J2MID_GHb_BEG1_input[2]),
	.A3 (J2MID_GHb_BEG1_input[3]),
	.S0 (ConfigBits[208+0]),
	.S0N (ConfigBits_N[208+0]),
	.S1 (ConfigBits[208+1]),
	.S1N (ConfigBits_N[208+1]),
	.X (J2MID_GHb_BEG1)
	);

// switch matrix multiplexer  J2MID_GHb_BEG2 		MUX-4
	assign J2MID_GHb_BEG2_input = {W2MID5,S2MID5,E2MID5,N2MID5};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_GHb_BEG2 (
	.A0 (J2MID_GHb_BEG2_input[0]),
	.A1 (J2MID_GHb_BEG2_input[1]),
	.A2 (J2MID_GHb_BEG2_input[2]),
	.A3 (J2MID_GHb_BEG2_input[3]),
	.S0 (ConfigBits[210+0]),
	.S0N (ConfigBits_N[210+0]),
	.S1 (ConfigBits[210+1]),
	.S1N (ConfigBits_N[210+1]),
	.X (J2MID_GHb_BEG2)
	);

// switch matrix multiplexer  J2MID_GHb_BEG3 		MUX-4
	assign J2MID_GHb_BEG3_input = {W2MID1,S2MID1,E2MID1,N2MID1};
	cus_mux41_buf inst_cus_mux41_buf_J2MID_GHb_BEG3 (
	.A0 (J2MID_GHb_BEG3_input[0]),
	.A1 (J2MID_GHb_BEG3_input[1]),
	.A2 (J2MID_GHb_BEG3_input[2]),
	.A3 (J2MID_GHb_BEG3_input[3]),
	.S0 (ConfigBits[212+0]),
	.S0N (ConfigBits_N[212+0]),
	.S1 (ConfigBits[212+1]),
	.S1N (ConfigBits_N[212+1]),
	.X (J2MID_GHb_BEG3)
	);

// switch matrix multiplexer  J2END_AB_BEG0 		MUX-4
	assign J2END_AB_BEG0_input = {W2END6,SS4END3,E2END6,N2END6};
	cus_mux41_buf inst_cus_mux41_buf_J2END_AB_BEG0 (
	.A0 (J2END_AB_BEG0_input[0]),
	.A1 (J2END_AB_BEG0_input[1]),
	.A2 (J2END_AB_BEG0_input[2]),
	.A3 (J2END_AB_BEG0_input[3]),
	.S0 (ConfigBits[214+0]),
	.S0N (ConfigBits_N[214+0]),
	.S1 (ConfigBits[214+1]),
	.S1N (ConfigBits_N[214+1]),
	.X (J2END_AB_BEG0)
	);

// switch matrix multiplexer  J2END_AB_BEG1 		MUX-4
	assign J2END_AB_BEG1_input = {W2END2,S2END2,E2END2,NN4END0};
	cus_mux41_buf inst_cus_mux41_buf_J2END_AB_BEG1 (
	.A0 (J2END_AB_BEG1_input[0]),
	.A1 (J2END_AB_BEG1_input[1]),
	.A2 (J2END_AB_BEG1_input[2]),
	.A3 (J2END_AB_BEG1_input[3]),
	.S0 (ConfigBits[216+0]),
	.S0N (ConfigBits_N[216+0]),
	.S1 (ConfigBits[216+1]),
	.S1N (ConfigBits_N[216+1]),
	.X (J2END_AB_BEG1)
	);

// switch matrix multiplexer  J2END_AB_BEG2 		MUX-4
	assign J2END_AB_BEG2_input = {W2END4,S2END4,EE4END0,N2END4};
	cus_mux41_buf inst_cus_mux41_buf_J2END_AB_BEG2 (
	.A0 (J2END_AB_BEG2_input[0]),
	.A1 (J2END_AB_BEG2_input[1]),
	.A2 (J2END_AB_BEG2_input[2]),
	.A3 (J2END_AB_BEG2_input[3]),
	.S0 (ConfigBits[218+0]),
	.S0N (ConfigBits_N[218+0]),
	.S1 (ConfigBits[218+1]),
	.S1N (ConfigBits_N[218+1]),
	.X (J2END_AB_BEG2)
	);

// switch matrix multiplexer  J2END_AB_BEG3 		MUX-4
	assign J2END_AB_BEG3_input = {WW4END3,S2END0,E2END0,N2END0};
	cus_mux41_buf inst_cus_mux41_buf_J2END_AB_BEG3 (
	.A0 (J2END_AB_BEG3_input[0]),
	.A1 (J2END_AB_BEG3_input[1]),
	.A2 (J2END_AB_BEG3_input[2]),
	.A3 (J2END_AB_BEG3_input[3]),
	.S0 (ConfigBits[220+0]),
	.S0N (ConfigBits_N[220+0]),
	.S1 (ConfigBits[220+1]),
	.S1N (ConfigBits_N[220+1]),
	.X (J2END_AB_BEG3)
	);

// switch matrix multiplexer  J2END_CD_BEG0 		MUX-4
	assign J2END_CD_BEG0_input = {W2END6,S2END6,E2END6,NN4END3};
	cus_mux41_buf inst_cus_mux41_buf_J2END_CD_BEG0 (
	.A0 (J2END_CD_BEG0_input[0]),
	.A1 (J2END_CD_BEG0_input[1]),
	.A2 (J2END_CD_BEG0_input[2]),
	.A3 (J2END_CD_BEG0_input[3]),
	.S0 (ConfigBits[222+0]),
	.S0N (ConfigBits_N[222+0]),
	.S1 (ConfigBits[222+1]),
	.S1N (ConfigBits_N[222+1]),
	.X (J2END_CD_BEG0)
	);

// switch matrix multiplexer  J2END_CD_BEG1 		MUX-4
	assign J2END_CD_BEG1_input = {WW4END2,S2END2,E2END2,N2END2};
	cus_mux41_buf inst_cus_mux41_buf_J2END_CD_BEG1 (
	.A0 (J2END_CD_BEG1_input[0]),
	.A1 (J2END_CD_BEG1_input[1]),
	.A2 (J2END_CD_BEG1_input[2]),
	.A3 (J2END_CD_BEG1_input[3]),
	.S0 (ConfigBits[224+0]),
	.S0N (ConfigBits_N[224+0]),
	.S1 (ConfigBits[224+1]),
	.S1N (ConfigBits_N[224+1]),
	.X (J2END_CD_BEG1)
	);

// switch matrix multiplexer  J2END_CD_BEG2 		MUX-4
	assign J2END_CD_BEG2_input = {W2END4,SS4END2,E2END4,N2END4};
	cus_mux41_buf inst_cus_mux41_buf_J2END_CD_BEG2 (
	.A0 (J2END_CD_BEG2_input[0]),
	.A1 (J2END_CD_BEG2_input[1]),
	.A2 (J2END_CD_BEG2_input[2]),
	.A3 (J2END_CD_BEG2_input[3]),
	.S0 (ConfigBits[226+0]),
	.S0N (ConfigBits_N[226+0]),
	.S1 (ConfigBits[226+1]),
	.S1N (ConfigBits_N[226+1]),
	.X (J2END_CD_BEG2)
	);

// switch matrix multiplexer  J2END_CD_BEG3 		MUX-4
	assign J2END_CD_BEG3_input = {W2END0,S2END0,EE4END1,N2END0};
	cus_mux41_buf inst_cus_mux41_buf_J2END_CD_BEG3 (
	.A0 (J2END_CD_BEG3_input[0]),
	.A1 (J2END_CD_BEG3_input[1]),
	.A2 (J2END_CD_BEG3_input[2]),
	.A3 (J2END_CD_BEG3_input[3]),
	.S0 (ConfigBits[228+0]),
	.S0N (ConfigBits_N[228+0]),
	.S1 (ConfigBits[228+1]),
	.S1N (ConfigBits_N[228+1]),
	.X (J2END_CD_BEG3)
	);

// switch matrix multiplexer  J2END_EF_BEG0 		MUX-4
	assign J2END_EF_BEG0_input = {W2END7,S2END7,EE4END2,N2END7};
	cus_mux41_buf inst_cus_mux41_buf_J2END_EF_BEG0 (
	.A0 (J2END_EF_BEG0_input[0]),
	.A1 (J2END_EF_BEG0_input[1]),
	.A2 (J2END_EF_BEG0_input[2]),
	.A3 (J2END_EF_BEG0_input[3]),
	.S0 (ConfigBits[230+0]),
	.S0N (ConfigBits_N[230+0]),
	.S1 (ConfigBits[230+1]),
	.S1N (ConfigBits_N[230+1]),
	.X (J2END_EF_BEG0)
	);

// switch matrix multiplexer  J2END_EF_BEG1 		MUX-4
	assign J2END_EF_BEG1_input = {WW4END1,S2END3,E2END3,N2END3};
	cus_mux41_buf inst_cus_mux41_buf_J2END_EF_BEG1 (
	.A0 (J2END_EF_BEG1_input[0]),
	.A1 (J2END_EF_BEG1_input[1]),
	.A2 (J2END_EF_BEG1_input[2]),
	.A3 (J2END_EF_BEG1_input[3]),
	.S0 (ConfigBits[232+0]),
	.S0N (ConfigBits_N[232+0]),
	.S1 (ConfigBits[232+1]),
	.S1N (ConfigBits_N[232+1]),
	.X (J2END_EF_BEG1)
	);

// switch matrix multiplexer  J2END_EF_BEG2 		MUX-4
	assign J2END_EF_BEG2_input = {W2END5,SS4END1,E2END5,N2END5};
	cus_mux41_buf inst_cus_mux41_buf_J2END_EF_BEG2 (
	.A0 (J2END_EF_BEG2_input[0]),
	.A1 (J2END_EF_BEG2_input[1]),
	.A2 (J2END_EF_BEG2_input[2]),
	.A3 (J2END_EF_BEG2_input[3]),
	.S0 (ConfigBits[234+0]),
	.S0N (ConfigBits_N[234+0]),
	.S1 (ConfigBits[234+1]),
	.S1N (ConfigBits_N[234+1]),
	.X (J2END_EF_BEG2)
	);

// switch matrix multiplexer  J2END_EF_BEG3 		MUX-4
	assign J2END_EF_BEG3_input = {W2END1,S2END1,E2END1,NN4END2};
	cus_mux41_buf inst_cus_mux41_buf_J2END_EF_BEG3 (
	.A0 (J2END_EF_BEG3_input[0]),
	.A1 (J2END_EF_BEG3_input[1]),
	.A2 (J2END_EF_BEG3_input[2]),
	.A3 (J2END_EF_BEG3_input[3]),
	.S0 (ConfigBits[236+0]),
	.S0N (ConfigBits_N[236+0]),
	.S1 (ConfigBits[236+1]),
	.S1N (ConfigBits_N[236+1]),
	.X (J2END_EF_BEG3)
	);

// switch matrix multiplexer  J2END_GH_BEG0 		MUX-4
	assign J2END_GH_BEG0_input = {WW4END0,S2END7,E2END7,N2END7};
	cus_mux41_buf inst_cus_mux41_buf_J2END_GH_BEG0 (
	.A0 (J2END_GH_BEG0_input[0]),
	.A1 (J2END_GH_BEG0_input[1]),
	.A2 (J2END_GH_BEG0_input[2]),
	.A3 (J2END_GH_BEG0_input[3]),
	.S0 (ConfigBits[238+0]),
	.S0N (ConfigBits_N[238+0]),
	.S1 (ConfigBits[238+1]),
	.S1N (ConfigBits_N[238+1]),
	.X (J2END_GH_BEG0)
	);

// switch matrix multiplexer  J2END_GH_BEG1 		MUX-4
	assign J2END_GH_BEG1_input = {W2END3,SS4END0,E2END3,N2END3};
	cus_mux41_buf inst_cus_mux41_buf_J2END_GH_BEG1 (
	.A0 (J2END_GH_BEG1_input[0]),
	.A1 (J2END_GH_BEG1_input[1]),
	.A2 (J2END_GH_BEG1_input[2]),
	.A3 (J2END_GH_BEG1_input[3]),
	.S0 (ConfigBits[240+0]),
	.S0N (ConfigBits_N[240+0]),
	.S1 (ConfigBits[240+1]),
	.S1N (ConfigBits_N[240+1]),
	.X (J2END_GH_BEG1)
	);

// switch matrix multiplexer  J2END_GH_BEG2 		MUX-4
	assign J2END_GH_BEG2_input = {W2END5,S2END5,E2END5,NN4END1};
	cus_mux41_buf inst_cus_mux41_buf_J2END_GH_BEG2 (
	.A0 (J2END_GH_BEG2_input[0]),
	.A1 (J2END_GH_BEG2_input[1]),
	.A2 (J2END_GH_BEG2_input[2]),
	.A3 (J2END_GH_BEG2_input[3]),
	.S0 (ConfigBits[242+0]),
	.S0N (ConfigBits_N[242+0]),
	.S1 (ConfigBits[242+1]),
	.S1N (ConfigBits_N[242+1]),
	.X (J2END_GH_BEG2)
	);

// switch matrix multiplexer  J2END_GH_BEG3 		MUX-4
	assign J2END_GH_BEG3_input = {W2END1,S2END1,EE4END3,N2END1};
	cus_mux41_buf inst_cus_mux41_buf_J2END_GH_BEG3 (
	.A0 (J2END_GH_BEG3_input[0]),
	.A1 (J2END_GH_BEG3_input[1]),
	.A2 (J2END_GH_BEG3_input[2]),
	.A3 (J2END_GH_BEG3_input[3]),
	.S0 (ConfigBits[244+0]),
	.S0N (ConfigBits_N[244+0]),
	.S1 (ConfigBits[244+1]),
	.S1N (ConfigBits_N[244+1]),
	.X (J2END_GH_BEG3)
	);

// switch matrix multiplexer  JN2BEG0 		MUX-16
	assign JN2BEG0_input = {W6END1,W2END1,SS4END1,E6END1,E2END1,E1END3,bot2top9,bot2top7,bot2top6,bot2top5,bot2top4,bot2top3,bot2top2,bot2top1,N4END1,N2END1};
	cus_mux161_buf inst_cus_mux161_buf_JN2BEG0 (
	.A0 (JN2BEG0_input[0]),
	.A1 (JN2BEG0_input[1]),
	.A2 (JN2BEG0_input[2]),
	.A3 (JN2BEG0_input[3]),
	.A4 (JN2BEG0_input[4]),
	.A5 (JN2BEG0_input[5]),
	.A6 (JN2BEG0_input[6]),
	.A7 (JN2BEG0_input[7]),
	.A8 (JN2BEG0_input[8]),
	.A9 (JN2BEG0_input[9]),
	.A10 (JN2BEG0_input[10]),
	.A11 (JN2BEG0_input[11]),
	.A12 (JN2BEG0_input[12]),
	.A13 (JN2BEG0_input[13]),
	.A14 (JN2BEG0_input[14]),
	.A15 (JN2BEG0_input[15]),
	.S0 (ConfigBits[246+0]),
	.S0N (ConfigBits_N[246+0]),
	.S1 (ConfigBits[246+1]),
	.S1N (ConfigBits_N[246+1]),
	.S2 (ConfigBits[246+2]),
	.S2N (ConfigBits_N[246+2]),
	.S3 (ConfigBits[246+3]),
	.S3N (ConfigBits_N[246+3]),
	.X (JN2BEG0)
	);

// switch matrix multiplexer  JN2BEG1 		MUX-16
	assign JN2BEG1_input = {W6END0,W2END2,S2END2,E6END0,E2END2,E1END0,bot2top8,bot2top7,bot2top6,bot2top5,bot2top4,bot2top3,bot2top2,bot2top0,N4END2,N2END2};
	cus_mux161_buf inst_cus_mux161_buf_JN2BEG1 (
	.A0 (JN2BEG1_input[0]),
	.A1 (JN2BEG1_input[1]),
	.A2 (JN2BEG1_input[2]),
	.A3 (JN2BEG1_input[3]),
	.A4 (JN2BEG1_input[4]),
	.A5 (JN2BEG1_input[5]),
	.A6 (JN2BEG1_input[6]),
	.A7 (JN2BEG1_input[7]),
	.A8 (JN2BEG1_input[8]),
	.A9 (JN2BEG1_input[9]),
	.A10 (JN2BEG1_input[10]),
	.A11 (JN2BEG1_input[11]),
	.A12 (JN2BEG1_input[12]),
	.A13 (JN2BEG1_input[13]),
	.A14 (JN2BEG1_input[14]),
	.A15 (JN2BEG1_input[15]),
	.S0 (ConfigBits[250+0]),
	.S0N (ConfigBits_N[250+0]),
	.S1 (ConfigBits[250+1]),
	.S1N (ConfigBits_N[250+1]),
	.S2 (ConfigBits[250+2]),
	.S2N (ConfigBits_N[250+2]),
	.S3 (ConfigBits[250+3]),
	.S3N (ConfigBits_N[250+3]),
	.X (JN2BEG1)
	);

// switch matrix multiplexer  JN2BEG2 		MUX-16
	assign JN2BEG2_input = {WW4END1,W2END3,S2END3,E6END1,E2END3,E1END1,bot2top9,bot2top7,bot2top6,bot2top5,bot2top4,bot2top3,bot2top1,bot2top0,N4END3,N2END3};
	cus_mux161_buf inst_cus_mux161_buf_JN2BEG2 (
	.A0 (JN2BEG2_input[0]),
	.A1 (JN2BEG2_input[1]),
	.A2 (JN2BEG2_input[2]),
	.A3 (JN2BEG2_input[3]),
	.A4 (JN2BEG2_input[4]),
	.A5 (JN2BEG2_input[5]),
	.A6 (JN2BEG2_input[6]),
	.A7 (JN2BEG2_input[7]),
	.A8 (JN2BEG2_input[8]),
	.A9 (JN2BEG2_input[9]),
	.A10 (JN2BEG2_input[10]),
	.A11 (JN2BEG2_input[11]),
	.A12 (JN2BEG2_input[12]),
	.A13 (JN2BEG2_input[13]),
	.A14 (JN2BEG2_input[14]),
	.A15 (JN2BEG2_input[15]),
	.S0 (ConfigBits[254+0]),
	.S0N (ConfigBits_N[254+0]),
	.S1 (ConfigBits[254+1]),
	.S1N (ConfigBits_N[254+1]),
	.S2 (ConfigBits[254+2]),
	.S2N (ConfigBits_N[254+2]),
	.S3 (ConfigBits[254+3]),
	.S3N (ConfigBits_N[254+3]),
	.X (JN2BEG2)
	);

// switch matrix multiplexer  JN2BEG3 		MUX-16
	assign JN2BEG3_input = {W6END0,W2END4,S2END4,E6END0,E2END4,E1END2,bot2top8,bot2top7,bot2top6,bot2top5,bot2top4,bot2top2,bot2top1,bot2top0,N4END0,N2END4};
	cus_mux161_buf inst_cus_mux161_buf_JN2BEG3 (
	.A0 (JN2BEG3_input[0]),
	.A1 (JN2BEG3_input[1]),
	.A2 (JN2BEG3_input[2]),
	.A3 (JN2BEG3_input[3]),
	.A4 (JN2BEG3_input[4]),
	.A5 (JN2BEG3_input[5]),
	.A6 (JN2BEG3_input[6]),
	.A7 (JN2BEG3_input[7]),
	.A8 (JN2BEG3_input[8]),
	.A9 (JN2BEG3_input[9]),
	.A10 (JN2BEG3_input[10]),
	.A11 (JN2BEG3_input[11]),
	.A12 (JN2BEG3_input[12]),
	.A13 (JN2BEG3_input[13]),
	.A14 (JN2BEG3_input[14]),
	.A15 (JN2BEG3_input[15]),
	.S0 (ConfigBits[258+0]),
	.S0N (ConfigBits_N[258+0]),
	.S1 (ConfigBits[258+1]),
	.S1N (ConfigBits_N[258+1]),
	.S2 (ConfigBits[258+2]),
	.S2N (ConfigBits_N[258+2]),
	.S3 (ConfigBits[258+3]),
	.S3N (ConfigBits_N[258+3]),
	.X (JN2BEG3)
	);

// switch matrix multiplexer  JN2BEG4 		MUX-16
	assign JN2BEG4_input = {W1END3,W1END1,S2END5,S1END1,E2END5,E1END1,bot2top9,bot2top7,bot2top6,bot2top5,bot2top3,bot2top2,bot2top1,bot2top0,N2END5,N1END1};
	cus_mux161_buf inst_cus_mux161_buf_JN2BEG4 (
	.A0 (JN2BEG4_input[0]),
	.A1 (JN2BEG4_input[1]),
	.A2 (JN2BEG4_input[2]),
	.A3 (JN2BEG4_input[3]),
	.A4 (JN2BEG4_input[4]),
	.A5 (JN2BEG4_input[5]),
	.A6 (JN2BEG4_input[6]),
	.A7 (JN2BEG4_input[7]),
	.A8 (JN2BEG4_input[8]),
	.A9 (JN2BEG4_input[9]),
	.A10 (JN2BEG4_input[10]),
	.A11 (JN2BEG4_input[11]),
	.A12 (JN2BEG4_input[12]),
	.A13 (JN2BEG4_input[13]),
	.A14 (JN2BEG4_input[14]),
	.A15 (JN2BEG4_input[15]),
	.S0 (ConfigBits[262+0]),
	.S0N (ConfigBits_N[262+0]),
	.S1 (ConfigBits[262+1]),
	.S1N (ConfigBits_N[262+1]),
	.S2 (ConfigBits[262+2]),
	.S2N (ConfigBits_N[262+2]),
	.S3 (ConfigBits[262+3]),
	.S3N (ConfigBits_N[262+3]),
	.X (JN2BEG4)
	);

// switch matrix multiplexer  JN2BEG5 		MUX-16
	assign JN2BEG5_input = {W1END2,W1END0,S2END6,S1END2,E2END6,E1END2,bot2top8,bot2top7,bot2top6,bot2top4,bot2top3,bot2top2,bot2top1,bot2top0,N2END6,N1END2};
	cus_mux161_buf inst_cus_mux161_buf_JN2BEG5 (
	.A0 (JN2BEG5_input[0]),
	.A1 (JN2BEG5_input[1]),
	.A2 (JN2BEG5_input[2]),
	.A3 (JN2BEG5_input[3]),
	.A4 (JN2BEG5_input[4]),
	.A5 (JN2BEG5_input[5]),
	.A6 (JN2BEG5_input[6]),
	.A7 (JN2BEG5_input[7]),
	.A8 (JN2BEG5_input[8]),
	.A9 (JN2BEG5_input[9]),
	.A10 (JN2BEG5_input[10]),
	.A11 (JN2BEG5_input[11]),
	.A12 (JN2BEG5_input[12]),
	.A13 (JN2BEG5_input[13]),
	.A14 (JN2BEG5_input[14]),
	.A15 (JN2BEG5_input[15]),
	.S0 (ConfigBits[266+0]),
	.S0N (ConfigBits_N[266+0]),
	.S1 (ConfigBits[266+1]),
	.S1N (ConfigBits_N[266+1]),
	.S2 (ConfigBits[266+2]),
	.S2N (ConfigBits_N[266+2]),
	.S3 (ConfigBits[266+3]),
	.S3N (ConfigBits_N[266+3]),
	.X (JN2BEG5)
	);

// switch matrix multiplexer  JN2BEG6 		MUX-16
	assign JN2BEG6_input = {W1END3,W1END1,S2END7,S1END3,E2END7,E1END3,bot2top9,bot2top7,bot2top5,bot2top4,bot2top3,bot2top2,bot2top1,bot2top0,N2END7,N1END3};
	cus_mux161_buf inst_cus_mux161_buf_JN2BEG6 (
	.A0 (JN2BEG6_input[0]),
	.A1 (JN2BEG6_input[1]),
	.A2 (JN2BEG6_input[2]),
	.A3 (JN2BEG6_input[3]),
	.A4 (JN2BEG6_input[4]),
	.A5 (JN2BEG6_input[5]),
	.A6 (JN2BEG6_input[6]),
	.A7 (JN2BEG6_input[7]),
	.A8 (JN2BEG6_input[8]),
	.A9 (JN2BEG6_input[9]),
	.A10 (JN2BEG6_input[10]),
	.A11 (JN2BEG6_input[11]),
	.A12 (JN2BEG6_input[12]),
	.A13 (JN2BEG6_input[13]),
	.A14 (JN2BEG6_input[14]),
	.A15 (JN2BEG6_input[15]),
	.S0 (ConfigBits[270+0]),
	.S0N (ConfigBits_N[270+0]),
	.S1 (ConfigBits[270+1]),
	.S1N (ConfigBits_N[270+1]),
	.S2 (ConfigBits[270+2]),
	.S2N (ConfigBits_N[270+2]),
	.S3 (ConfigBits[270+3]),
	.S3N (ConfigBits_N[270+3]),
	.X (JN2BEG6)
	);

// switch matrix multiplexer  JN2BEG7 		MUX-16
	assign JN2BEG7_input = {W1END2,W1END0,S2END0,S1END0,EE4END0,E1END0,bot2top8,bot2top6,bot2top5,bot2top4,bot2top3,bot2top2,bot2top1,bot2top0,N2END0,N1END0};
	cus_mux161_buf inst_cus_mux161_buf_JN2BEG7 (
	.A0 (JN2BEG7_input[0]),
	.A1 (JN2BEG7_input[1]),
	.A2 (JN2BEG7_input[2]),
	.A3 (JN2BEG7_input[3]),
	.A4 (JN2BEG7_input[4]),
	.A5 (JN2BEG7_input[5]),
	.A6 (JN2BEG7_input[6]),
	.A7 (JN2BEG7_input[7]),
	.A8 (JN2BEG7_input[8]),
	.A9 (JN2BEG7_input[9]),
	.A10 (JN2BEG7_input[10]),
	.A11 (JN2BEG7_input[11]),
	.A12 (JN2BEG7_input[12]),
	.A13 (JN2BEG7_input[13]),
	.A14 (JN2BEG7_input[14]),
	.A15 (JN2BEG7_input[15]),
	.S0 (ConfigBits[274+0]),
	.S0N (ConfigBits_N[274+0]),
	.S1 (ConfigBits[274+1]),
	.S1N (ConfigBits_N[274+1]),
	.S2 (ConfigBits[274+2]),
	.S2N (ConfigBits_N[274+2]),
	.S3 (ConfigBits[274+3]),
	.S3N (ConfigBits_N[274+3]),
	.X (JN2BEG7)
	);

// switch matrix multiplexer  JE2BEG0 		MUX-16
	assign JE2BEG0_input = {W6END1,W2END1,S2END1,E6END1,EE4END1,bot2top8,bot2top7,bot2top6,bot2top5,bot2top4,bot2top3,bot2top2,bot2top1,N4END1,N2END1,N1END3};
	cus_mux161_buf inst_cus_mux161_buf_JE2BEG0 (
	.A0 (JE2BEG0_input[0]),
	.A1 (JE2BEG0_input[1]),
	.A2 (JE2BEG0_input[2]),
	.A3 (JE2BEG0_input[3]),
	.A4 (JE2BEG0_input[4]),
	.A5 (JE2BEG0_input[5]),
	.A6 (JE2BEG0_input[6]),
	.A7 (JE2BEG0_input[7]),
	.A8 (JE2BEG0_input[8]),
	.A9 (JE2BEG0_input[9]),
	.A10 (JE2BEG0_input[10]),
	.A11 (JE2BEG0_input[11]),
	.A12 (JE2BEG0_input[12]),
	.A13 (JE2BEG0_input[13]),
	.A14 (JE2BEG0_input[14]),
	.A15 (JE2BEG0_input[15]),
	.S0 (ConfigBits[278+0]),
	.S0N (ConfigBits_N[278+0]),
	.S1 (ConfigBits[278+1]),
	.S1N (ConfigBits_N[278+1]),
	.S2 (ConfigBits[278+2]),
	.S2N (ConfigBits_N[278+2]),
	.S3 (ConfigBits[278+3]),
	.S3N (ConfigBits_N[278+3]),
	.X (JE2BEG0)
	);

// switch matrix multiplexer  JE2BEG1 		MUX-16
	assign JE2BEG1_input = {WW4END3,W2END2,S2END2,E6END0,E2END2,bot2top9,bot2top7,bot2top6,bot2top5,bot2top4,bot2top3,bot2top2,bot2top0,N4END2,N2END2,N1END0};
	cus_mux161_buf inst_cus_mux161_buf_JE2BEG1 (
	.A0 (JE2BEG1_input[0]),
	.A1 (JE2BEG1_input[1]),
	.A2 (JE2BEG1_input[2]),
	.A3 (JE2BEG1_input[3]),
	.A4 (JE2BEG1_input[4]),
	.A5 (JE2BEG1_input[5]),
	.A6 (JE2BEG1_input[6]),
	.A7 (JE2BEG1_input[7]),
	.A8 (JE2BEG1_input[8]),
	.A9 (JE2BEG1_input[9]),
	.A10 (JE2BEG1_input[10]),
	.A11 (JE2BEG1_input[11]),
	.A12 (JE2BEG1_input[12]),
	.A13 (JE2BEG1_input[13]),
	.A14 (JE2BEG1_input[14]),
	.A15 (JE2BEG1_input[15]),
	.S0 (ConfigBits[282+0]),
	.S0N (ConfigBits_N[282+0]),
	.S1 (ConfigBits[282+1]),
	.S1N (ConfigBits_N[282+1]),
	.S2 (ConfigBits[282+2]),
	.S2N (ConfigBits_N[282+2]),
	.S3 (ConfigBits[282+3]),
	.S3N (ConfigBits_N[282+3]),
	.X (JE2BEG1)
	);

// switch matrix multiplexer  JE2BEG2 		MUX-16
	assign JE2BEG2_input = {W6END1,W2END3,S2END3,E6END1,E2END3,bot2top8,bot2top7,bot2top6,bot2top5,bot2top4,bot2top3,bot2top1,bot2top0,N4END3,N2END3,N1END1};
	cus_mux161_buf inst_cus_mux161_buf_JE2BEG2 (
	.A0 (JE2BEG2_input[0]),
	.A1 (JE2BEG2_input[1]),
	.A2 (JE2BEG2_input[2]),
	.A3 (JE2BEG2_input[3]),
	.A4 (JE2BEG2_input[4]),
	.A5 (JE2BEG2_input[5]),
	.A6 (JE2BEG2_input[6]),
	.A7 (JE2BEG2_input[7]),
	.A8 (JE2BEG2_input[8]),
	.A9 (JE2BEG2_input[9]),
	.A10 (JE2BEG2_input[10]),
	.A11 (JE2BEG2_input[11]),
	.A12 (JE2BEG2_input[12]),
	.A13 (JE2BEG2_input[13]),
	.A14 (JE2BEG2_input[14]),
	.A15 (JE2BEG2_input[15]),
	.S0 (ConfigBits[286+0]),
	.S0N (ConfigBits_N[286+0]),
	.S1 (ConfigBits[286+1]),
	.S1N (ConfigBits_N[286+1]),
	.S2 (ConfigBits[286+2]),
	.S2N (ConfigBits_N[286+2]),
	.S3 (ConfigBits[286+3]),
	.S3N (ConfigBits_N[286+3]),
	.X (JE2BEG2)
	);

// switch matrix multiplexer  JE2BEG3 		MUX-16
	assign JE2BEG3_input = {W6END0,W2END4,S2END4,E6END0,E2END4,bot2top9,bot2top7,bot2top6,bot2top5,bot2top4,bot2top2,bot2top1,bot2top0,N4END0,N2END4,N1END2};
	cus_mux161_buf inst_cus_mux161_buf_JE2BEG3 (
	.A0 (JE2BEG3_input[0]),
	.A1 (JE2BEG3_input[1]),
	.A2 (JE2BEG3_input[2]),
	.A3 (JE2BEG3_input[3]),
	.A4 (JE2BEG3_input[4]),
	.A5 (JE2BEG3_input[5]),
	.A6 (JE2BEG3_input[6]),
	.A7 (JE2BEG3_input[7]),
	.A8 (JE2BEG3_input[8]),
	.A9 (JE2BEG3_input[9]),
	.A10 (JE2BEG3_input[10]),
	.A11 (JE2BEG3_input[11]),
	.A12 (JE2BEG3_input[12]),
	.A13 (JE2BEG3_input[13]),
	.A14 (JE2BEG3_input[14]),
	.A15 (JE2BEG3_input[15]),
	.S0 (ConfigBits[290+0]),
	.S0N (ConfigBits_N[290+0]),
	.S1 (ConfigBits[290+1]),
	.S1N (ConfigBits_N[290+1]),
	.S2 (ConfigBits[290+2]),
	.S2N (ConfigBits_N[290+2]),
	.S3 (ConfigBits[290+3]),
	.S3N (ConfigBits_N[290+3]),
	.X (JE2BEG3)
	);

// switch matrix multiplexer  JE2BEG4 		MUX-16
	assign JE2BEG4_input = {W1END1,S2END5,S1END3,S1END1,E2END5,E1END1,bot2top8,bot2top7,bot2top6,bot2top5,bot2top3,bot2top2,bot2top1,bot2top0,N2END5,N1END1};
	cus_mux161_buf inst_cus_mux161_buf_JE2BEG4 (
	.A0 (JE2BEG4_input[0]),
	.A1 (JE2BEG4_input[1]),
	.A2 (JE2BEG4_input[2]),
	.A3 (JE2BEG4_input[3]),
	.A4 (JE2BEG4_input[4]),
	.A5 (JE2BEG4_input[5]),
	.A6 (JE2BEG4_input[6]),
	.A7 (JE2BEG4_input[7]),
	.A8 (JE2BEG4_input[8]),
	.A9 (JE2BEG4_input[9]),
	.A10 (JE2BEG4_input[10]),
	.A11 (JE2BEG4_input[11]),
	.A12 (JE2BEG4_input[12]),
	.A13 (JE2BEG4_input[13]),
	.A14 (JE2BEG4_input[14]),
	.A15 (JE2BEG4_input[15]),
	.S0 (ConfigBits[294+0]),
	.S0N (ConfigBits_N[294+0]),
	.S1 (ConfigBits[294+1]),
	.S1N (ConfigBits_N[294+1]),
	.S2 (ConfigBits[294+2]),
	.S2N (ConfigBits_N[294+2]),
	.S3 (ConfigBits[294+3]),
	.S3N (ConfigBits_N[294+3]),
	.X (JE2BEG4)
	);

// switch matrix multiplexer  JE2BEG5 		MUX-16
	assign JE2BEG5_input = {W1END2,S2END6,S1END2,S1END0,E2END6,E1END2,bot2top9,bot2top7,bot2top6,bot2top4,bot2top3,bot2top2,bot2top1,bot2top0,N2END6,N1END2};
	cus_mux161_buf inst_cus_mux161_buf_JE2BEG5 (
	.A0 (JE2BEG5_input[0]),
	.A1 (JE2BEG5_input[1]),
	.A2 (JE2BEG5_input[2]),
	.A3 (JE2BEG5_input[3]),
	.A4 (JE2BEG5_input[4]),
	.A5 (JE2BEG5_input[5]),
	.A6 (JE2BEG5_input[6]),
	.A7 (JE2BEG5_input[7]),
	.A8 (JE2BEG5_input[8]),
	.A9 (JE2BEG5_input[9]),
	.A10 (JE2BEG5_input[10]),
	.A11 (JE2BEG5_input[11]),
	.A12 (JE2BEG5_input[12]),
	.A13 (JE2BEG5_input[13]),
	.A14 (JE2BEG5_input[14]),
	.A15 (JE2BEG5_input[15]),
	.S0 (ConfigBits[298+0]),
	.S0N (ConfigBits_N[298+0]),
	.S1 (ConfigBits[298+1]),
	.S1N (ConfigBits_N[298+1]),
	.S2 (ConfigBits[298+2]),
	.S2N (ConfigBits_N[298+2]),
	.S3 (ConfigBits[298+3]),
	.S3N (ConfigBits_N[298+3]),
	.X (JE2BEG5)
	);

// switch matrix multiplexer  JE2BEG6 		MUX-16
	assign JE2BEG6_input = {W1END3,S2END7,S1END3,S1END1,E2END7,E1END3,bot2top8,bot2top7,bot2top5,bot2top4,bot2top3,bot2top2,bot2top1,bot2top0,N2END7,N1END3};
	cus_mux161_buf inst_cus_mux161_buf_JE2BEG6 (
	.A0 (JE2BEG6_input[0]),
	.A1 (JE2BEG6_input[1]),
	.A2 (JE2BEG6_input[2]),
	.A3 (JE2BEG6_input[3]),
	.A4 (JE2BEG6_input[4]),
	.A5 (JE2BEG6_input[5]),
	.A6 (JE2BEG6_input[6]),
	.A7 (JE2BEG6_input[7]),
	.A8 (JE2BEG6_input[8]),
	.A9 (JE2BEG6_input[9]),
	.A10 (JE2BEG6_input[10]),
	.A11 (JE2BEG6_input[11]),
	.A12 (JE2BEG6_input[12]),
	.A13 (JE2BEG6_input[13]),
	.A14 (JE2BEG6_input[14]),
	.A15 (JE2BEG6_input[15]),
	.S0 (ConfigBits[302+0]),
	.S0N (ConfigBits_N[302+0]),
	.S1 (ConfigBits[302+1]),
	.S1N (ConfigBits_N[302+1]),
	.S2 (ConfigBits[302+2]),
	.S2N (ConfigBits_N[302+2]),
	.S3 (ConfigBits[302+3]),
	.S3N (ConfigBits_N[302+3]),
	.X (JE2BEG6)
	);

// switch matrix multiplexer  JE2BEG7 		MUX-16
	assign JE2BEG7_input = {WW4END0,SS4END0,S1END2,S1END0,E2END0,E1END0,bot2top9,bot2top6,bot2top5,bot2top4,bot2top3,bot2top2,bot2top1,bot2top0,N2END0,N1END0};
	cus_mux161_buf inst_cus_mux161_buf_JE2BEG7 (
	.A0 (JE2BEG7_input[0]),
	.A1 (JE2BEG7_input[1]),
	.A2 (JE2BEG7_input[2]),
	.A3 (JE2BEG7_input[3]),
	.A4 (JE2BEG7_input[4]),
	.A5 (JE2BEG7_input[5]),
	.A6 (JE2BEG7_input[6]),
	.A7 (JE2BEG7_input[7]),
	.A8 (JE2BEG7_input[8]),
	.A9 (JE2BEG7_input[9]),
	.A10 (JE2BEG7_input[10]),
	.A11 (JE2BEG7_input[11]),
	.A12 (JE2BEG7_input[12]),
	.A13 (JE2BEG7_input[13]),
	.A14 (JE2BEG7_input[14]),
	.A15 (JE2BEG7_input[15]),
	.S0 (ConfigBits[306+0]),
	.S0N (ConfigBits_N[306+0]),
	.S1 (ConfigBits[306+1]),
	.S1N (ConfigBits_N[306+1]),
	.S2 (ConfigBits[306+2]),
	.S2N (ConfigBits_N[306+2]),
	.S3 (ConfigBits[306+3]),
	.S3N (ConfigBits_N[306+3]),
	.X (JE2BEG7)
	);

// switch matrix multiplexer  JS2BEG0 		MUX-16
	assign JS2BEG0_input = {W6END1,W2END1,S4END1,S2END1,E6END1,E2END1,E1END3,bot2top9,bot2top7,bot2top6,bot2top5,bot2top4,bot2top3,bot2top2,bot2top1,NN4END1};
	cus_mux161_buf inst_cus_mux161_buf_JS2BEG0 (
	.A0 (JS2BEG0_input[0]),
	.A1 (JS2BEG0_input[1]),
	.A2 (JS2BEG0_input[2]),
	.A3 (JS2BEG0_input[3]),
	.A4 (JS2BEG0_input[4]),
	.A5 (JS2BEG0_input[5]),
	.A6 (JS2BEG0_input[6]),
	.A7 (JS2BEG0_input[7]),
	.A8 (JS2BEG0_input[8]),
	.A9 (JS2BEG0_input[9]),
	.A10 (JS2BEG0_input[10]),
	.A11 (JS2BEG0_input[11]),
	.A12 (JS2BEG0_input[12]),
	.A13 (JS2BEG0_input[13]),
	.A14 (JS2BEG0_input[14]),
	.A15 (JS2BEG0_input[15]),
	.S0 (ConfigBits[310+0]),
	.S0N (ConfigBits_N[310+0]),
	.S1 (ConfigBits[310+1]),
	.S1N (ConfigBits_N[310+1]),
	.S2 (ConfigBits[310+2]),
	.S2N (ConfigBits_N[310+2]),
	.S3 (ConfigBits[310+3]),
	.S3N (ConfigBits_N[310+3]),
	.X (JS2BEG0)
	);

// switch matrix multiplexer  JS2BEG1 		MUX-16
	assign JS2BEG1_input = {W6END0,W2END2,SS4END2,S4END2,E6END0,EE4END2,E1END0,bot2top8,bot2top7,bot2top6,bot2top5,bot2top4,bot2top3,bot2top2,bot2top0,NN4END2};
	cus_mux161_buf inst_cus_mux161_buf_JS2BEG1 (
	.A0 (JS2BEG1_input[0]),
	.A1 (JS2BEG1_input[1]),
	.A2 (JS2BEG1_input[2]),
	.A3 (JS2BEG1_input[3]),
	.A4 (JS2BEG1_input[4]),
	.A5 (JS2BEG1_input[5]),
	.A6 (JS2BEG1_input[6]),
	.A7 (JS2BEG1_input[7]),
	.A8 (JS2BEG1_input[8]),
	.A9 (JS2BEG1_input[9]),
	.A10 (JS2BEG1_input[10]),
	.A11 (JS2BEG1_input[11]),
	.A12 (JS2BEG1_input[12]),
	.A13 (JS2BEG1_input[13]),
	.A14 (JS2BEG1_input[14]),
	.A15 (JS2BEG1_input[15]),
	.S0 (ConfigBits[314+0]),
	.S0N (ConfigBits_N[314+0]),
	.S1 (ConfigBits[314+1]),
	.S1N (ConfigBits_N[314+1]),
	.S2 (ConfigBits[314+2]),
	.S2N (ConfigBits_N[314+2]),
	.S3 (ConfigBits[314+3]),
	.S3N (ConfigBits_N[314+3]),
	.X (JS2BEG1)
	);

// switch matrix multiplexer  JS2BEG2 		MUX-16
	assign JS2BEG2_input = {W6END1,W2END3,S4END3,S2END3,E6END1,E2END3,E1END1,bot2top9,bot2top7,bot2top6,bot2top5,bot2top4,bot2top3,bot2top1,bot2top0,NN4END3};
	cus_mux161_buf inst_cus_mux161_buf_JS2BEG2 (
	.A0 (JS2BEG2_input[0]),
	.A1 (JS2BEG2_input[1]),
	.A2 (JS2BEG2_input[2]),
	.A3 (JS2BEG2_input[3]),
	.A4 (JS2BEG2_input[4]),
	.A5 (JS2BEG2_input[5]),
	.A6 (JS2BEG2_input[6]),
	.A7 (JS2BEG2_input[7]),
	.A8 (JS2BEG2_input[8]),
	.A9 (JS2BEG2_input[9]),
	.A10 (JS2BEG2_input[10]),
	.A11 (JS2BEG2_input[11]),
	.A12 (JS2BEG2_input[12]),
	.A13 (JS2BEG2_input[13]),
	.A14 (JS2BEG2_input[14]),
	.A15 (JS2BEG2_input[15]),
	.S0 (ConfigBits[318+0]),
	.S0N (ConfigBits_N[318+0]),
	.S1 (ConfigBits[318+1]),
	.S1N (ConfigBits_N[318+1]),
	.S2 (ConfigBits[318+2]),
	.S2N (ConfigBits_N[318+2]),
	.S3 (ConfigBits[318+3]),
	.S3N (ConfigBits_N[318+3]),
	.X (JS2BEG2)
	);

// switch matrix multiplexer  JS2BEG3 		MUX-16
	assign JS2BEG3_input = {WW4END2,W2END4,S4END0,S2END4,E6END0,E2END4,E1END2,bot2top8,bot2top7,bot2top6,bot2top5,bot2top4,bot2top2,bot2top1,bot2top0,N2END4};
	cus_mux161_buf inst_cus_mux161_buf_JS2BEG3 (
	.A0 (JS2BEG3_input[0]),
	.A1 (JS2BEG3_input[1]),
	.A2 (JS2BEG3_input[2]),
	.A3 (JS2BEG3_input[3]),
	.A4 (JS2BEG3_input[4]),
	.A5 (JS2BEG3_input[5]),
	.A6 (JS2BEG3_input[6]),
	.A7 (JS2BEG3_input[7]),
	.A8 (JS2BEG3_input[8]),
	.A9 (JS2BEG3_input[9]),
	.A10 (JS2BEG3_input[10]),
	.A11 (JS2BEG3_input[11]),
	.A12 (JS2BEG3_input[12]),
	.A13 (JS2BEG3_input[13]),
	.A14 (JS2BEG3_input[14]),
	.A15 (JS2BEG3_input[15]),
	.S0 (ConfigBits[322+0]),
	.S0N (ConfigBits_N[322+0]),
	.S1 (ConfigBits[322+1]),
	.S1N (ConfigBits_N[322+1]),
	.S2 (ConfigBits[322+2]),
	.S2N (ConfigBits_N[322+2]),
	.S3 (ConfigBits[322+3]),
	.S3N (ConfigBits_N[322+3]),
	.X (JS2BEG3)
	);

// switch matrix multiplexer  JS2BEG4 		MUX-16
	assign JS2BEG4_input = {W1END3,W1END1,S2END5,S1END1,E2END5,E1END1,bot2top9,bot2top7,bot2top6,bot2top5,bot2top3,bot2top2,bot2top1,bot2top0,N2END5,N1END1};
	cus_mux161_buf inst_cus_mux161_buf_JS2BEG4 (
	.A0 (JS2BEG4_input[0]),
	.A1 (JS2BEG4_input[1]),
	.A2 (JS2BEG4_input[2]),
	.A3 (JS2BEG4_input[3]),
	.A4 (JS2BEG4_input[4]),
	.A5 (JS2BEG4_input[5]),
	.A6 (JS2BEG4_input[6]),
	.A7 (JS2BEG4_input[7]),
	.A8 (JS2BEG4_input[8]),
	.A9 (JS2BEG4_input[9]),
	.A10 (JS2BEG4_input[10]),
	.A11 (JS2BEG4_input[11]),
	.A12 (JS2BEG4_input[12]),
	.A13 (JS2BEG4_input[13]),
	.A14 (JS2BEG4_input[14]),
	.A15 (JS2BEG4_input[15]),
	.S0 (ConfigBits[326+0]),
	.S0N (ConfigBits_N[326+0]),
	.S1 (ConfigBits[326+1]),
	.S1N (ConfigBits_N[326+1]),
	.S2 (ConfigBits[326+2]),
	.S2N (ConfigBits_N[326+2]),
	.S3 (ConfigBits[326+3]),
	.S3N (ConfigBits_N[326+3]),
	.X (JS2BEG4)
	);

// switch matrix multiplexer  JS2BEG5 		MUX-16
	assign JS2BEG5_input = {W1END2,W1END0,S2END6,S1END2,E2END6,E1END2,bot2top8,bot2top7,bot2top6,bot2top4,bot2top3,bot2top2,bot2top1,bot2top0,N2END6,N1END2};
	cus_mux161_buf inst_cus_mux161_buf_JS2BEG5 (
	.A0 (JS2BEG5_input[0]),
	.A1 (JS2BEG5_input[1]),
	.A2 (JS2BEG5_input[2]),
	.A3 (JS2BEG5_input[3]),
	.A4 (JS2BEG5_input[4]),
	.A5 (JS2BEG5_input[5]),
	.A6 (JS2BEG5_input[6]),
	.A7 (JS2BEG5_input[7]),
	.A8 (JS2BEG5_input[8]),
	.A9 (JS2BEG5_input[9]),
	.A10 (JS2BEG5_input[10]),
	.A11 (JS2BEG5_input[11]),
	.A12 (JS2BEG5_input[12]),
	.A13 (JS2BEG5_input[13]),
	.A14 (JS2BEG5_input[14]),
	.A15 (JS2BEG5_input[15]),
	.S0 (ConfigBits[330+0]),
	.S0N (ConfigBits_N[330+0]),
	.S1 (ConfigBits[330+1]),
	.S1N (ConfigBits_N[330+1]),
	.S2 (ConfigBits[330+2]),
	.S2N (ConfigBits_N[330+2]),
	.S3 (ConfigBits[330+3]),
	.S3N (ConfigBits_N[330+3]),
	.X (JS2BEG5)
	);

// switch matrix multiplexer  JS2BEG6 		MUX-16
	assign JS2BEG6_input = {W1END3,W1END1,S2END7,S1END3,E2END7,E1END3,bot2top9,bot2top7,bot2top5,bot2top4,bot2top3,bot2top2,bot2top1,bot2top0,N2END7,N1END3};
	cus_mux161_buf inst_cus_mux161_buf_JS2BEG6 (
	.A0 (JS2BEG6_input[0]),
	.A1 (JS2BEG6_input[1]),
	.A2 (JS2BEG6_input[2]),
	.A3 (JS2BEG6_input[3]),
	.A4 (JS2BEG6_input[4]),
	.A5 (JS2BEG6_input[5]),
	.A6 (JS2BEG6_input[6]),
	.A7 (JS2BEG6_input[7]),
	.A8 (JS2BEG6_input[8]),
	.A9 (JS2BEG6_input[9]),
	.A10 (JS2BEG6_input[10]),
	.A11 (JS2BEG6_input[11]),
	.A12 (JS2BEG6_input[12]),
	.A13 (JS2BEG6_input[13]),
	.A14 (JS2BEG6_input[14]),
	.A15 (JS2BEG6_input[15]),
	.S0 (ConfigBits[334+0]),
	.S0N (ConfigBits_N[334+0]),
	.S1 (ConfigBits[334+1]),
	.S1N (ConfigBits_N[334+1]),
	.S2 (ConfigBits[334+2]),
	.S2N (ConfigBits_N[334+2]),
	.S3 (ConfigBits[334+3]),
	.S3N (ConfigBits_N[334+3]),
	.X (JS2BEG6)
	);

// switch matrix multiplexer  JS2BEG7 		MUX-16
	assign JS2BEG7_input = {W1END2,W1END0,S2END0,S1END0,E2END0,E1END0,bot2top8,bot2top6,bot2top5,bot2top4,bot2top3,bot2top2,bot2top1,bot2top0,N2END0,N1END0};
	cus_mux161_buf inst_cus_mux161_buf_JS2BEG7 (
	.A0 (JS2BEG7_input[0]),
	.A1 (JS2BEG7_input[1]),
	.A2 (JS2BEG7_input[2]),
	.A3 (JS2BEG7_input[3]),
	.A4 (JS2BEG7_input[4]),
	.A5 (JS2BEG7_input[5]),
	.A6 (JS2BEG7_input[6]),
	.A7 (JS2BEG7_input[7]),
	.A8 (JS2BEG7_input[8]),
	.A9 (JS2BEG7_input[9]),
	.A10 (JS2BEG7_input[10]),
	.A11 (JS2BEG7_input[11]),
	.A12 (JS2BEG7_input[12]),
	.A13 (JS2BEG7_input[13]),
	.A14 (JS2BEG7_input[14]),
	.A15 (JS2BEG7_input[15]),
	.S0 (ConfigBits[338+0]),
	.S0N (ConfigBits_N[338+0]),
	.S1 (ConfigBits[338+1]),
	.S1N (ConfigBits_N[338+1]),
	.S2 (ConfigBits[338+2]),
	.S2N (ConfigBits_N[338+2]),
	.S3 (ConfigBits[338+3]),
	.S3N (ConfigBits_N[338+3]),
	.X (JS2BEG7)
	);

// switch matrix multiplexer  JW2BEG0 		MUX-16
	assign JW2BEG0_input = {W6END1,W2END1,S4END1,S2END1,E6END1,E2END1,bot2top8,bot2top7,bot2top6,bot2top5,bot2top4,bot2top3,bot2top2,bot2top1,N2END1,N1END3};
	cus_mux161_buf inst_cus_mux161_buf_JW2BEG0 (
	.A0 (JW2BEG0_input[0]),
	.A1 (JW2BEG0_input[1]),
	.A2 (JW2BEG0_input[2]),
	.A3 (JW2BEG0_input[3]),
	.A4 (JW2BEG0_input[4]),
	.A5 (JW2BEG0_input[5]),
	.A6 (JW2BEG0_input[6]),
	.A7 (JW2BEG0_input[7]),
	.A8 (JW2BEG0_input[8]),
	.A9 (JW2BEG0_input[9]),
	.A10 (JW2BEG0_input[10]),
	.A11 (JW2BEG0_input[11]),
	.A12 (JW2BEG0_input[12]),
	.A13 (JW2BEG0_input[13]),
	.A14 (JW2BEG0_input[14]),
	.A15 (JW2BEG0_input[15]),
	.S0 (ConfigBits[342+0]),
	.S0N (ConfigBits_N[342+0]),
	.S1 (ConfigBits[342+1]),
	.S1N (ConfigBits_N[342+1]),
	.S2 (ConfigBits[342+2]),
	.S2N (ConfigBits_N[342+2]),
	.S3 (ConfigBits[342+3]),
	.S3N (ConfigBits_N[342+3]),
	.X (JW2BEG0)
	);

// switch matrix multiplexer  JW2BEG1 		MUX-16
	assign JW2BEG1_input = {W6END0,W2END2,S4END2,S2END2,E6END0,E2END2,bot2top9,bot2top7,bot2top6,bot2top5,bot2top4,bot2top3,bot2top2,bot2top0,N2END2,N1END0};
	cus_mux161_buf inst_cus_mux161_buf_JW2BEG1 (
	.A0 (JW2BEG1_input[0]),
	.A1 (JW2BEG1_input[1]),
	.A2 (JW2BEG1_input[2]),
	.A3 (JW2BEG1_input[3]),
	.A4 (JW2BEG1_input[4]),
	.A5 (JW2BEG1_input[5]),
	.A6 (JW2BEG1_input[6]),
	.A7 (JW2BEG1_input[7]),
	.A8 (JW2BEG1_input[8]),
	.A9 (JW2BEG1_input[9]),
	.A10 (JW2BEG1_input[10]),
	.A11 (JW2BEG1_input[11]),
	.A12 (JW2BEG1_input[12]),
	.A13 (JW2BEG1_input[13]),
	.A14 (JW2BEG1_input[14]),
	.A15 (JW2BEG1_input[15]),
	.S0 (ConfigBits[346+0]),
	.S0N (ConfigBits_N[346+0]),
	.S1 (ConfigBits[346+1]),
	.S1N (ConfigBits_N[346+1]),
	.S2 (ConfigBits[346+2]),
	.S2N (ConfigBits_N[346+2]),
	.S3 (ConfigBits[346+3]),
	.S3N (ConfigBits_N[346+3]),
	.X (JW2BEG1)
	);

// switch matrix multiplexer  JW2BEG2 		MUX-16
	assign JW2BEG2_input = {W6END1,W2END3,S4END3,S2END3,E6END1,E2END3,bot2top8,bot2top7,bot2top6,bot2top5,bot2top4,bot2top3,bot2top1,bot2top0,N2END3,N1END1};
	cus_mux161_buf inst_cus_mux161_buf_JW2BEG2 (
	.A0 (JW2BEG2_input[0]),
	.A1 (JW2BEG2_input[1]),
	.A2 (JW2BEG2_input[2]),
	.A3 (JW2BEG2_input[3]),
	.A4 (JW2BEG2_input[4]),
	.A5 (JW2BEG2_input[5]),
	.A6 (JW2BEG2_input[6]),
	.A7 (JW2BEG2_input[7]),
	.A8 (JW2BEG2_input[8]),
	.A9 (JW2BEG2_input[9]),
	.A10 (JW2BEG2_input[10]),
	.A11 (JW2BEG2_input[11]),
	.A12 (JW2BEG2_input[12]),
	.A13 (JW2BEG2_input[13]),
	.A14 (JW2BEG2_input[14]),
	.A15 (JW2BEG2_input[15]),
	.S0 (ConfigBits[350+0]),
	.S0N (ConfigBits_N[350+0]),
	.S1 (ConfigBits[350+1]),
	.S1N (ConfigBits_N[350+1]),
	.S2 (ConfigBits[350+2]),
	.S2N (ConfigBits_N[350+2]),
	.S3 (ConfigBits[350+3]),
	.S3N (ConfigBits_N[350+3]),
	.X (JW2BEG2)
	);

// switch matrix multiplexer  JW2BEG3 		MUX-16
	assign JW2BEG3_input = {W6END0,W2END4,S4END0,S2END4,E6END0,E2END4,bot2top9,bot2top7,bot2top6,bot2top5,bot2top4,bot2top2,bot2top1,bot2top0,N2END4,N1END2};
	cus_mux161_buf inst_cus_mux161_buf_JW2BEG3 (
	.A0 (JW2BEG3_input[0]),
	.A1 (JW2BEG3_input[1]),
	.A2 (JW2BEG3_input[2]),
	.A3 (JW2BEG3_input[3]),
	.A4 (JW2BEG3_input[4]),
	.A5 (JW2BEG3_input[5]),
	.A6 (JW2BEG3_input[6]),
	.A7 (JW2BEG3_input[7]),
	.A8 (JW2BEG3_input[8]),
	.A9 (JW2BEG3_input[9]),
	.A10 (JW2BEG3_input[10]),
	.A11 (JW2BEG3_input[11]),
	.A12 (JW2BEG3_input[12]),
	.A13 (JW2BEG3_input[13]),
	.A14 (JW2BEG3_input[14]),
	.A15 (JW2BEG3_input[15]),
	.S0 (ConfigBits[354+0]),
	.S0N (ConfigBits_N[354+0]),
	.S1 (ConfigBits[354+1]),
	.S1N (ConfigBits_N[354+1]),
	.S2 (ConfigBits[354+2]),
	.S2N (ConfigBits_N[354+2]),
	.S3 (ConfigBits[354+3]),
	.S3N (ConfigBits_N[354+3]),
	.X (JW2BEG3)
	);

// switch matrix multiplexer  JW2BEG4 		MUX-16
	assign JW2BEG4_input = {W1END1,S2END5,S1END3,S1END1,E2END5,E1END1,bot2top8,bot2top7,bot2top6,bot2top5,bot2top3,bot2top2,bot2top1,bot2top0,N2END5,N1END1};
	cus_mux161_buf inst_cus_mux161_buf_JW2BEG4 (
	.A0 (JW2BEG4_input[0]),
	.A1 (JW2BEG4_input[1]),
	.A2 (JW2BEG4_input[2]),
	.A3 (JW2BEG4_input[3]),
	.A4 (JW2BEG4_input[4]),
	.A5 (JW2BEG4_input[5]),
	.A6 (JW2BEG4_input[6]),
	.A7 (JW2BEG4_input[7]),
	.A8 (JW2BEG4_input[8]),
	.A9 (JW2BEG4_input[9]),
	.A10 (JW2BEG4_input[10]),
	.A11 (JW2BEG4_input[11]),
	.A12 (JW2BEG4_input[12]),
	.A13 (JW2BEG4_input[13]),
	.A14 (JW2BEG4_input[14]),
	.A15 (JW2BEG4_input[15]),
	.S0 (ConfigBits[358+0]),
	.S0N (ConfigBits_N[358+0]),
	.S1 (ConfigBits[358+1]),
	.S1N (ConfigBits_N[358+1]),
	.S2 (ConfigBits[358+2]),
	.S2N (ConfigBits_N[358+2]),
	.S3 (ConfigBits[358+3]),
	.S3N (ConfigBits_N[358+3]),
	.X (JW2BEG4)
	);

// switch matrix multiplexer  JW2BEG5 		MUX-16
	assign JW2BEG5_input = {W1END2,S2END6,S1END2,S1END0,E2END6,E1END2,bot2top9,bot2top7,bot2top6,bot2top4,bot2top3,bot2top2,bot2top1,bot2top0,N2END6,N1END2};
	cus_mux161_buf inst_cus_mux161_buf_JW2BEG5 (
	.A0 (JW2BEG5_input[0]),
	.A1 (JW2BEG5_input[1]),
	.A2 (JW2BEG5_input[2]),
	.A3 (JW2BEG5_input[3]),
	.A4 (JW2BEG5_input[4]),
	.A5 (JW2BEG5_input[5]),
	.A6 (JW2BEG5_input[6]),
	.A7 (JW2BEG5_input[7]),
	.A8 (JW2BEG5_input[8]),
	.A9 (JW2BEG5_input[9]),
	.A10 (JW2BEG5_input[10]),
	.A11 (JW2BEG5_input[11]),
	.A12 (JW2BEG5_input[12]),
	.A13 (JW2BEG5_input[13]),
	.A14 (JW2BEG5_input[14]),
	.A15 (JW2BEG5_input[15]),
	.S0 (ConfigBits[362+0]),
	.S0N (ConfigBits_N[362+0]),
	.S1 (ConfigBits[362+1]),
	.S1N (ConfigBits_N[362+1]),
	.S2 (ConfigBits[362+2]),
	.S2N (ConfigBits_N[362+2]),
	.S3 (ConfigBits[362+3]),
	.S3N (ConfigBits_N[362+3]),
	.X (JW2BEG5)
	);

// switch matrix multiplexer  JW2BEG6 		MUX-16
	assign JW2BEG6_input = {W1END3,S2END7,S1END3,S1END1,E2END7,E1END3,bot2top8,bot2top7,bot2top5,bot2top4,bot2top3,bot2top2,bot2top1,bot2top0,N2END7,N1END3};
	cus_mux161_buf inst_cus_mux161_buf_JW2BEG6 (
	.A0 (JW2BEG6_input[0]),
	.A1 (JW2BEG6_input[1]),
	.A2 (JW2BEG6_input[2]),
	.A3 (JW2BEG6_input[3]),
	.A4 (JW2BEG6_input[4]),
	.A5 (JW2BEG6_input[5]),
	.A6 (JW2BEG6_input[6]),
	.A7 (JW2BEG6_input[7]),
	.A8 (JW2BEG6_input[8]),
	.A9 (JW2BEG6_input[9]),
	.A10 (JW2BEG6_input[10]),
	.A11 (JW2BEG6_input[11]),
	.A12 (JW2BEG6_input[12]),
	.A13 (JW2BEG6_input[13]),
	.A14 (JW2BEG6_input[14]),
	.A15 (JW2BEG6_input[15]),
	.S0 (ConfigBits[366+0]),
	.S0N (ConfigBits_N[366+0]),
	.S1 (ConfigBits[366+1]),
	.S1N (ConfigBits_N[366+1]),
	.S2 (ConfigBits[366+2]),
	.S2N (ConfigBits_N[366+2]),
	.S3 (ConfigBits[366+3]),
	.S3N (ConfigBits_N[366+3]),
	.X (JW2BEG6)
	);

// switch matrix multiplexer  JW2BEG7 		MUX-16
	assign JW2BEG7_input = {W1END0,S2END0,S1END2,S1END0,E2END0,E1END0,bot2top9,bot2top6,bot2top5,bot2top4,bot2top3,bot2top2,bot2top1,bot2top0,N2END0,N1END0};
	cus_mux161_buf inst_cus_mux161_buf_JW2BEG7 (
	.A0 (JW2BEG7_input[0]),
	.A1 (JW2BEG7_input[1]),
	.A2 (JW2BEG7_input[2]),
	.A3 (JW2BEG7_input[3]),
	.A4 (JW2BEG7_input[4]),
	.A5 (JW2BEG7_input[5]),
	.A6 (JW2BEG7_input[6]),
	.A7 (JW2BEG7_input[7]),
	.A8 (JW2BEG7_input[8]),
	.A9 (JW2BEG7_input[9]),
	.A10 (JW2BEG7_input[10]),
	.A11 (JW2BEG7_input[11]),
	.A12 (JW2BEG7_input[12]),
	.A13 (JW2BEG7_input[13]),
	.A14 (JW2BEG7_input[14]),
	.A15 (JW2BEG7_input[15]),
	.S0 (ConfigBits[370+0]),
	.S0N (ConfigBits_N[370+0]),
	.S1 (ConfigBits[370+1]),
	.S1N (ConfigBits_N[370+1]),
	.S2 (ConfigBits[370+2]),
	.S2N (ConfigBits_N[370+2]),
	.S3 (ConfigBits[370+3]),
	.S3N (ConfigBits_N[370+3]),
	.X (JW2BEG7)
	);

// switch matrix multiplexer  J_l_AB_BEG0 		MUX-4
	assign J_l_AB_BEG0_input = {JN2END1,WW4END0,S4END3,NN4END3};
	cus_mux41_buf inst_cus_mux41_buf_J_l_AB_BEG0 (
	.A0 (J_l_AB_BEG0_input[0]),
	.A1 (J_l_AB_BEG0_input[1]),
	.A2 (J_l_AB_BEG0_input[2]),
	.A3 (J_l_AB_BEG0_input[3]),
	.S0 (ConfigBits[374+0]),
	.S0N (ConfigBits_N[374+0]),
	.S1 (ConfigBits[374+1]),
	.S1N (ConfigBits_N[374+1]),
	.X (J_l_AB_BEG0)
	);

// switch matrix multiplexer  J_l_AB_BEG1 		MUX-4
	assign J_l_AB_BEG1_input = {JE2END1,W2END7,S4END2,EE4END2};
	cus_mux41_buf inst_cus_mux41_buf_J_l_AB_BEG1 (
	.A0 (J_l_AB_BEG1_input[0]),
	.A1 (J_l_AB_BEG1_input[1]),
	.A2 (J_l_AB_BEG1_input[2]),
	.A3 (J_l_AB_BEG1_input[3]),
	.S0 (ConfigBits[376+0]),
	.S0N (ConfigBits_N[376+0]),
	.S1 (ConfigBits[376+1]),
	.S1N (ConfigBits_N[376+1]),
	.X (J_l_AB_BEG1)
	);

// switch matrix multiplexer  J_l_AB_BEG2 		MUX-4
	assign J_l_AB_BEG2_input = {JS2END1,W6END1,E6END1,N4END1};
	cus_mux41_buf inst_cus_mux41_buf_J_l_AB_BEG2 (
	.A0 (J_l_AB_BEG2_input[0]),
	.A1 (J_l_AB_BEG2_input[1]),
	.A2 (J_l_AB_BEG2_input[2]),
	.A3 (J_l_AB_BEG2_input[3]),
	.S0 (ConfigBits[378+0]),
	.S0N (ConfigBits_N[378+0]),
	.S1 (ConfigBits[378+1]),
	.S1N (ConfigBits_N[378+1]),
	.X (J_l_AB_BEG2)
	);

// switch matrix multiplexer  J_l_AB_BEG3 		MUX-4
	assign J_l_AB_BEG3_input = {JW2END1,S4END0,E6END0,N4END0};
	cus_mux41_buf inst_cus_mux41_buf_J_l_AB_BEG3 (
	.A0 (J_l_AB_BEG3_input[0]),
	.A1 (J_l_AB_BEG3_input[1]),
	.A2 (J_l_AB_BEG3_input[2]),
	.A3 (J_l_AB_BEG3_input[3]),
	.S0 (ConfigBits[380+0]),
	.S0N (ConfigBits_N[380+0]),
	.S1 (ConfigBits[380+1]),
	.S1N (ConfigBits_N[380+1]),
	.X (J_l_AB_BEG3)
	);

// switch matrix multiplexer  J_l_CD_BEG0 		MUX-4
	assign J_l_CD_BEG0_input = {JN2END2,WW4END2,SS4END3,E2END3};
	cus_mux41_buf inst_cus_mux41_buf_J_l_CD_BEG0 (
	.A0 (J_l_CD_BEG0_input[0]),
	.A1 (J_l_CD_BEG0_input[1]),
	.A2 (J_l_CD_BEG0_input[2]),
	.A3 (J_l_CD_BEG0_input[3]),
	.S0 (ConfigBits[382+0]),
	.S0N (ConfigBits_N[382+0]),
	.S1 (ConfigBits[382+1]),
	.S1N (ConfigBits_N[382+1]),
	.X (J_l_CD_BEG0)
	);

// switch matrix multiplexer  J_l_CD_BEG1 		MUX-4
	assign J_l_CD_BEG1_input = {JE2END2,W2END7,E2END2,N4END2};
	cus_mux41_buf inst_cus_mux41_buf_J_l_CD_BEG1 (
	.A0 (J_l_CD_BEG1_input[0]),
	.A1 (J_l_CD_BEG1_input[1]),
	.A2 (J_l_CD_BEG1_input[2]),
	.A3 (J_l_CD_BEG1_input[3]),
	.S0 (ConfigBits[384+0]),
	.S0N (ConfigBits_N[384+0]),
	.S1 (ConfigBits[384+1]),
	.S1N (ConfigBits_N[384+1]),
	.X (J_l_CD_BEG1)
	);

// switch matrix multiplexer  J_l_CD_BEG2 		MUX-4
	assign J_l_CD_BEG2_input = {JS2END2,S4END1,EE4END1,NN4END1};
	cus_mux41_buf inst_cus_mux41_buf_J_l_CD_BEG2 (
	.A0 (J_l_CD_BEG2_input[0]),
	.A1 (J_l_CD_BEG2_input[1]),
	.A2 (J_l_CD_BEG2_input[2]),
	.A3 (J_l_CD_BEG2_input[3]),
	.S0 (ConfigBits[386+0]),
	.S0N (ConfigBits_N[386+0]),
	.S1 (ConfigBits[386+1]),
	.S1N (ConfigBits_N[386+1]),
	.X (J_l_CD_BEG2)
	);

// switch matrix multiplexer  J_l_CD_BEG3 		MUX-4
	assign J_l_CD_BEG3_input = {JW2END2,W6END0,SS4END0,N4END0};
	cus_mux41_buf inst_cus_mux41_buf_J_l_CD_BEG3 (
	.A0 (J_l_CD_BEG3_input[0]),
	.A1 (J_l_CD_BEG3_input[1]),
	.A2 (J_l_CD_BEG3_input[2]),
	.A3 (J_l_CD_BEG3_input[3]),
	.S0 (ConfigBits[388+0]),
	.S0N (ConfigBits_N[388+0]),
	.S1 (ConfigBits[388+1]),
	.S1N (ConfigBits_N[388+1]),
	.X (J_l_CD_BEG3)
	);

// switch matrix multiplexer  J_l_EF_BEG0 		MUX-4
	assign J_l_EF_BEG0_input = {JN2END3,W2END3,E2END3,N4END3};
	cus_mux41_buf inst_cus_mux41_buf_J_l_EF_BEG0 (
	.A0 (J_l_EF_BEG0_input[0]),
	.A1 (J_l_EF_BEG0_input[1]),
	.A2 (J_l_EF_BEG0_input[2]),
	.A3 (J_l_EF_BEG0_input[3]),
	.S0 (ConfigBits[390+0]),
	.S0N (ConfigBits_N[390+0]),
	.S1 (ConfigBits[390+1]),
	.S1N (ConfigBits_N[390+1]),
	.X (J_l_EF_BEG0)
	);

// switch matrix multiplexer  J_l_EF_BEG1 		MUX-4
	assign J_l_EF_BEG1_input = {JE2END3,S4END2,E2END2,NN4END2};
	cus_mux41_buf inst_cus_mux41_buf_J_l_EF_BEG1 (
	.A0 (J_l_EF_BEG1_input[0]),
	.A1 (J_l_EF_BEG1_input[1]),
	.A2 (J_l_EF_BEG1_input[2]),
	.A3 (J_l_EF_BEG1_input[3]),
	.S0 (ConfigBits[392+0]),
	.S0N (ConfigBits_N[392+0]),
	.S1 (ConfigBits[392+1]),
	.S1N (ConfigBits_N[392+1]),
	.X (J_l_EF_BEG1)
	);

// switch matrix multiplexer  J_l_EF_BEG2 		MUX-4
	assign J_l_EF_BEG2_input = {JS2END3,W2END4,SS4END1,N4END1};
	cus_mux41_buf inst_cus_mux41_buf_J_l_EF_BEG2 (
	.A0 (J_l_EF_BEG2_input[0]),
	.A1 (J_l_EF_BEG2_input[1]),
	.A2 (J_l_EF_BEG2_input[2]),
	.A3 (J_l_EF_BEG2_input[3]),
	.S0 (ConfigBits[394+0]),
	.S0N (ConfigBits_N[394+0]),
	.S1 (ConfigBits[394+1]),
	.S1N (ConfigBits_N[394+1]),
	.X (J_l_EF_BEG2)
	);

// switch matrix multiplexer  J_l_EF_BEG3 		MUX-4
	assign J_l_EF_BEG3_input = {JW2END3,WW4END1,S4END0,EE4END3};
	cus_mux41_buf inst_cus_mux41_buf_J_l_EF_BEG3 (
	.A0 (J_l_EF_BEG3_input[0]),
	.A1 (J_l_EF_BEG3_input[1]),
	.A2 (J_l_EF_BEG3_input[2]),
	.A3 (J_l_EF_BEG3_input[3]),
	.S0 (ConfigBits[396+0]),
	.S0N (ConfigBits_N[396+0]),
	.S1 (ConfigBits[396+1]),
	.S1N (ConfigBits_N[396+1]),
	.X (J_l_EF_BEG3)
	);

// switch matrix multiplexer  J_l_GH_BEG0 		MUX-4
	assign J_l_GH_BEG0_input = {JN2END4,S4END3,EE4END0,N4END3};
	cus_mux41_buf inst_cus_mux41_buf_J_l_GH_BEG0 (
	.A0 (J_l_GH_BEG0_input[0]),
	.A1 (J_l_GH_BEG0_input[1]),
	.A2 (J_l_GH_BEG0_input[2]),
	.A3 (J_l_GH_BEG0_input[3]),
	.S0 (ConfigBits[398+0]),
	.S0N (ConfigBits_N[398+0]),
	.S1 (ConfigBits[398+1]),
	.S1N (ConfigBits_N[398+1]),
	.X (J_l_GH_BEG0)
	);

// switch matrix multiplexer  J_l_GH_BEG1 		MUX-4
	assign J_l_GH_BEG1_input = {JE2END4,W2END2,SS4END2,N4END2};
	cus_mux41_buf inst_cus_mux41_buf_J_l_GH_BEG1 (
	.A0 (J_l_GH_BEG1_input[0]),
	.A1 (J_l_GH_BEG1_input[1]),
	.A2 (J_l_GH_BEG1_input[2]),
	.A3 (J_l_GH_BEG1_input[3]),
	.S0 (ConfigBits[400+0]),
	.S0N (ConfigBits_N[400+0]),
	.S1 (ConfigBits[400+1]),
	.S1N (ConfigBits_N[400+1]),
	.X (J_l_GH_BEG1)
	);

// switch matrix multiplexer  J_l_GH_BEG2 		MUX-4
	assign J_l_GH_BEG2_input = {JS2END4,WW4END3,S4END1,E6END1};
	cus_mux41_buf inst_cus_mux41_buf_J_l_GH_BEG2 (
	.A0 (J_l_GH_BEG2_input[0]),
	.A1 (J_l_GH_BEG2_input[1]),
	.A2 (J_l_GH_BEG2_input[2]),
	.A3 (J_l_GH_BEG2_input[3]),
	.S0 (ConfigBits[402+0]),
	.S0N (ConfigBits_N[402+0]),
	.S1 (ConfigBits[402+1]),
	.S1N (ConfigBits_N[402+1]),
	.X (J_l_GH_BEG2)
	);

// switch matrix multiplexer  J_l_GH_BEG3 		MUX-4
	assign J_l_GH_BEG3_input = {JW2END4,W2END0,E6END0,NN4END0};
	cus_mux41_buf inst_cus_mux41_buf_J_l_GH_BEG3 (
	.A0 (J_l_GH_BEG3_input[0]),
	.A1 (J_l_GH_BEG3_input[1]),
	.A2 (J_l_GH_BEG3_input[2]),
	.A3 (J_l_GH_BEG3_input[3]),
	.S0 (ConfigBits[404+0]),
	.S0N (ConfigBits_N[404+0]),
	.S1 (ConfigBits[404+1]),
	.S1N (ConfigBits_N[404+1]),
	.X (J_l_GH_BEG3)
	);

	assign DEBUG_select_N1BEG0 = ConfigBits[1:0];
	assign DEBUG_select_N1BEG1 = ConfigBits[3:2];
	assign DEBUG_select_N1BEG2 = ConfigBits[5:4];
	assign DEBUG_select_N1BEG3 = ConfigBits[7:6];
	assign DEBUG_select_N4BEG0 = ConfigBits[9:8];
	assign DEBUG_select_N4BEG1 = ConfigBits[11:10];
	assign DEBUG_select_N4BEG2 = ConfigBits[13:12];
	assign DEBUG_select_N4BEG3 = ConfigBits[15:14];
	assign DEBUG_select_NN4BEG0 = ConfigBits[18:16];
	assign DEBUG_select_NN4BEG1 = ConfigBits[21:19];
	assign DEBUG_select_NN4BEG2 = ConfigBits[24:22];
	assign DEBUG_select_NN4BEG3 = ConfigBits[27:25];
	assign DEBUG_select_E1BEG0 = ConfigBits[29:28];
	assign DEBUG_select_E1BEG1 = ConfigBits[31:30];
	assign DEBUG_select_E1BEG2 = ConfigBits[33:32];
	assign DEBUG_select_E1BEG3 = ConfigBits[35:34];
	assign DEBUG_select_EE4BEG0 = ConfigBits[38:36];
	assign DEBUG_select_EE4BEG1 = ConfigBits[41:39];
	assign DEBUG_select_EE4BEG2 = ConfigBits[44:42];
	assign DEBUG_select_EE4BEG3 = ConfigBits[47:45];
	assign DEBUG_select_E6BEG0 = ConfigBits[51:48];
	assign DEBUG_select_E6BEG1 = ConfigBits[55:52];
	assign DEBUG_select_S1BEG0 = ConfigBits[57:56];
	assign DEBUG_select_S1BEG1 = ConfigBits[59:58];
	assign DEBUG_select_S1BEG2 = ConfigBits[61:60];
	assign DEBUG_select_S1BEG3 = ConfigBits[63:62];
	assign DEBUG_select_S4BEG0 = ConfigBits[65:64];
	assign DEBUG_select_S4BEG1 = ConfigBits[67:66];
	assign DEBUG_select_S4BEG2 = ConfigBits[69:68];
	assign DEBUG_select_S4BEG3 = ConfigBits[71:70];
	assign DEBUG_select_SS4BEG0 = ConfigBits[74:72];
	assign DEBUG_select_SS4BEG1 = ConfigBits[77:75];
	assign DEBUG_select_SS4BEG2 = ConfigBits[80:78];
	assign DEBUG_select_SS4BEG3 = ConfigBits[83:81];
	assign DEBUG_select_top2bot0 = ConfigBits[85:84];
	assign DEBUG_select_top2bot1 = ConfigBits[87:86];
	assign DEBUG_select_top2bot2 = ConfigBits[89:88];
	assign DEBUG_select_top2bot3 = ConfigBits[91:90];
	assign DEBUG_select_top2bot4 = ConfigBits[93:92];
	assign DEBUG_select_top2bot5 = ConfigBits[95:94];
	assign DEBUG_select_top2bot6 = ConfigBits[97:96];
	assign DEBUG_select_top2bot7 = ConfigBits[99:98];
	assign DEBUG_select_top2bot8 = ConfigBits[101:100];
	assign DEBUG_select_top2bot9 = ConfigBits[103:102];
	assign DEBUG_select_top2bot10 = ConfigBits[105:104];
	assign DEBUG_select_top2bot11 = ConfigBits[107:106];
	assign DEBUG_select_top2bot12 = ConfigBits[109:108];
	assign DEBUG_select_top2bot13 = ConfigBits[111:110];
	assign DEBUG_select_top2bot14 = ConfigBits[113:112];
	assign DEBUG_select_top2bot15 = ConfigBits[115:114];
	assign DEBUG_select_top2bot16 = ConfigBits[118:116];
	assign DEBUG_select_top2bot17 = ConfigBits[121:119];
	assign DEBUG_select_W1BEG0 = ConfigBits[123:122];
	assign DEBUG_select_W1BEG1 = ConfigBits[125:124];
	assign DEBUG_select_W1BEG2 = ConfigBits[127:126];
	assign DEBUG_select_W1BEG3 = ConfigBits[129:128];
	assign DEBUG_select_WW4BEG0 = ConfigBits[132:130];
	assign DEBUG_select_WW4BEG1 = ConfigBits[135:133];
	assign DEBUG_select_WW4BEG2 = ConfigBits[138:136];
	assign DEBUG_select_WW4BEG3 = ConfigBits[141:139];
	assign DEBUG_select_W6BEG0 = ConfigBits[145:142];
	assign DEBUG_select_W6BEG1 = ConfigBits[149:146];
	assign DEBUG_select_J2MID_ABa_BEG0 = ConfigBits[151:150];
	assign DEBUG_select_J2MID_ABa_BEG1 = ConfigBits[153:152];
	assign DEBUG_select_J2MID_ABa_BEG2 = ConfigBits[155:154];
	assign DEBUG_select_J2MID_ABa_BEG3 = ConfigBits[157:156];
	assign DEBUG_select_J2MID_CDa_BEG0 = ConfigBits[159:158];
	assign DEBUG_select_J2MID_CDa_BEG1 = ConfigBits[161:160];
	assign DEBUG_select_J2MID_CDa_BEG2 = ConfigBits[163:162];
	assign DEBUG_select_J2MID_CDa_BEG3 = ConfigBits[165:164];
	assign DEBUG_select_J2MID_EFa_BEG0 = ConfigBits[167:166];
	assign DEBUG_select_J2MID_EFa_BEG1 = ConfigBits[169:168];
	assign DEBUG_select_J2MID_EFa_BEG2 = ConfigBits[171:170];
	assign DEBUG_select_J2MID_EFa_BEG3 = ConfigBits[173:172];
	assign DEBUG_select_J2MID_GHa_BEG0 = ConfigBits[175:174];
	assign DEBUG_select_J2MID_GHa_BEG1 = ConfigBits[177:176];
	assign DEBUG_select_J2MID_GHa_BEG2 = ConfigBits[179:178];
	assign DEBUG_select_J2MID_GHa_BEG3 = ConfigBits[181:180];
	assign DEBUG_select_J2MID_ABb_BEG0 = ConfigBits[183:182];
	assign DEBUG_select_J2MID_ABb_BEG1 = ConfigBits[185:184];
	assign DEBUG_select_J2MID_ABb_BEG2 = ConfigBits[187:186];
	assign DEBUG_select_J2MID_ABb_BEG3 = ConfigBits[189:188];
	assign DEBUG_select_J2MID_CDb_BEG0 = ConfigBits[191:190];
	assign DEBUG_select_J2MID_CDb_BEG1 = ConfigBits[193:192];
	assign DEBUG_select_J2MID_CDb_BEG2 = ConfigBits[195:194];
	assign DEBUG_select_J2MID_CDb_BEG3 = ConfigBits[197:196];
	assign DEBUG_select_J2MID_EFb_BEG0 = ConfigBits[199:198];
	assign DEBUG_select_J2MID_EFb_BEG1 = ConfigBits[201:200];
	assign DEBUG_select_J2MID_EFb_BEG2 = ConfigBits[203:202];
	assign DEBUG_select_J2MID_EFb_BEG3 = ConfigBits[205:204];
	assign DEBUG_select_J2MID_GHb_BEG0 = ConfigBits[207:206];
	assign DEBUG_select_J2MID_GHb_BEG1 = ConfigBits[209:208];
	assign DEBUG_select_J2MID_GHb_BEG2 = ConfigBits[211:210];
	assign DEBUG_select_J2MID_GHb_BEG3 = ConfigBits[213:212];
	assign DEBUG_select_J2END_AB_BEG0 = ConfigBits[215:214];
	assign DEBUG_select_J2END_AB_BEG1 = ConfigBits[217:216];
	assign DEBUG_select_J2END_AB_BEG2 = ConfigBits[219:218];
	assign DEBUG_select_J2END_AB_BEG3 = ConfigBits[221:220];
	assign DEBUG_select_J2END_CD_BEG0 = ConfigBits[223:222];
	assign DEBUG_select_J2END_CD_BEG1 = ConfigBits[225:224];
	assign DEBUG_select_J2END_CD_BEG2 = ConfigBits[227:226];
	assign DEBUG_select_J2END_CD_BEG3 = ConfigBits[229:228];
	assign DEBUG_select_J2END_EF_BEG0 = ConfigBits[231:230];
	assign DEBUG_select_J2END_EF_BEG1 = ConfigBits[233:232];
	assign DEBUG_select_J2END_EF_BEG2 = ConfigBits[235:234];
	assign DEBUG_select_J2END_EF_BEG3 = ConfigBits[237:236];
	assign DEBUG_select_J2END_GH_BEG0 = ConfigBits[239:238];
	assign DEBUG_select_J2END_GH_BEG1 = ConfigBits[241:240];
	assign DEBUG_select_J2END_GH_BEG2 = ConfigBits[243:242];
	assign DEBUG_select_J2END_GH_BEG3 = ConfigBits[245:244];
	assign DEBUG_select_JN2BEG0 = ConfigBits[249:246];
	assign DEBUG_select_JN2BEG1 = ConfigBits[253:250];
	assign DEBUG_select_JN2BEG2 = ConfigBits[257:254];
	assign DEBUG_select_JN2BEG3 = ConfigBits[261:258];
	assign DEBUG_select_JN2BEG4 = ConfigBits[265:262];
	assign DEBUG_select_JN2BEG5 = ConfigBits[269:266];
	assign DEBUG_select_JN2BEG6 = ConfigBits[273:270];
	assign DEBUG_select_JN2BEG7 = ConfigBits[277:274];
	assign DEBUG_select_JE2BEG0 = ConfigBits[281:278];
	assign DEBUG_select_JE2BEG1 = ConfigBits[285:282];
	assign DEBUG_select_JE2BEG2 = ConfigBits[289:286];
	assign DEBUG_select_JE2BEG3 = ConfigBits[293:290];
	assign DEBUG_select_JE2BEG4 = ConfigBits[297:294];
	assign DEBUG_select_JE2BEG5 = ConfigBits[301:298];
	assign DEBUG_select_JE2BEG6 = ConfigBits[305:302];
	assign DEBUG_select_JE2BEG7 = ConfigBits[309:306];
	assign DEBUG_select_JS2BEG0 = ConfigBits[313:310];
	assign DEBUG_select_JS2BEG1 = ConfigBits[317:314];
	assign DEBUG_select_JS2BEG2 = ConfigBits[321:318];
	assign DEBUG_select_JS2BEG3 = ConfigBits[325:322];
	assign DEBUG_select_JS2BEG4 = ConfigBits[329:326];
	assign DEBUG_select_JS2BEG5 = ConfigBits[333:330];
	assign DEBUG_select_JS2BEG6 = ConfigBits[337:334];
	assign DEBUG_select_JS2BEG7 = ConfigBits[341:338];
	assign DEBUG_select_JW2BEG0 = ConfigBits[345:342];
	assign DEBUG_select_JW2BEG1 = ConfigBits[349:346];
	assign DEBUG_select_JW2BEG2 = ConfigBits[353:350];
	assign DEBUG_select_JW2BEG3 = ConfigBits[357:354];
	assign DEBUG_select_JW2BEG4 = ConfigBits[361:358];
	assign DEBUG_select_JW2BEG5 = ConfigBits[365:362];
	assign DEBUG_select_JW2BEG6 = ConfigBits[369:366];
	assign DEBUG_select_JW2BEG7 = ConfigBits[373:370];
	assign DEBUG_select_J_l_AB_BEG0 = ConfigBits[375:374];
	assign DEBUG_select_J_l_AB_BEG1 = ConfigBits[377:376];
	assign DEBUG_select_J_l_AB_BEG2 = ConfigBits[379:378];
	assign DEBUG_select_J_l_AB_BEG3 = ConfigBits[381:380];
	assign DEBUG_select_J_l_CD_BEG0 = ConfigBits[383:382];
	assign DEBUG_select_J_l_CD_BEG1 = ConfigBits[385:384];
	assign DEBUG_select_J_l_CD_BEG2 = ConfigBits[387:386];
	assign DEBUG_select_J_l_CD_BEG3 = ConfigBits[389:388];
	assign DEBUG_select_J_l_EF_BEG0 = ConfigBits[391:390];
	assign DEBUG_select_J_l_EF_BEG1 = ConfigBits[393:392];
	assign DEBUG_select_J_l_EF_BEG2 = ConfigBits[395:394];
	assign DEBUG_select_J_l_EF_BEG3 = ConfigBits[397:396];
	assign DEBUG_select_J_l_GH_BEG0 = ConfigBits[399:398];
	assign DEBUG_select_J_l_GH_BEG1 = ConfigBits[401:400];
	assign DEBUG_select_J_l_GH_BEG2 = ConfigBits[403:402];
	assign DEBUG_select_J_l_GH_BEG3 = ConfigBits[405:404];

endmodule
