library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.my_package.all;

entity LUT4c_latch_config is
    -- Generic (LUT_SIZE : integer := 4);	
    Port (      -- IMPORTANT: this has to be in a dedicated line
	I0	: in	STD_LOGIC; -- LUT inputs
	I1	: in	STD_LOGIC;
	I2	: in	STD_LOGIC;
	I3	: in	STD_LOGIC;
	O	: out	STD_LOGIC; -- LUT output (combinatorial or FF)
	Ci	: in	STD_LOGIC; -- carry chain input
	Co	: out	STD_LOGIC; -- carry chain output
	UserCLK : in	STD_LOGIC; -- EXTERNAL -- the EXTERNAL keyword will send this signal all the way to top
	-- GLOBAL all primitive pins that are connected to the switch matrix have to go before the GLOBAL label
	MODE	: in 	 STD_LOGIC;	 -- 1 configuration, 0 action
	CONFin	: in 	 STD_LOGIC;
	CONFout	: out 	 STD_LOGIC;
	CLK	: in 	 STD_LOGIC
	);
end entity LUT4c_latch_config;

architecture Behavioral of LUT4c_latch_config is

constant LUT_SIZE : integer := 4; 
constant N_LUT_flops : integer := 2 ** LUT_SIZE; 


signal LUT_values : std_logic_vector(N_LUT_flops-1 downto 0);

signal LUT_index : unsigned(LUT_SIZE-1 downto 0);

signal LUT_out : std_logic;
signal LUT_flop  : std_logic;
signal I0mux              : std_logic;	-- normal input '0', or carry input '1'
signal c_out_mux, c_I0mux : std_logic;	-- extra configuration bits
signal ConfigBits :	 std_logic_vector( 16+2-1 downto 0 );
signal ConfigBitsInput :	 std_logic_vector( 16+2-1 downto 0 );

begin

-- The lookup tables are daisy-chained to a shift register made from latches

ConfigBitsInput <= ConfigBits(ConfigBits'high-1 downto 0) & CONFin; 

L: for k in 0 to 8 generate               
		inst_LHQD1a : LHQD1              
		Port Map(              
		D    => ConfigBitsInput(k*2),              
		E    => CLK,               
		Q    => ConfigBits(k*2) );                 
              
		inst_LHQD1b : LHQD1              
		Port Map(              
		D    => ConfigBitsInput((k*2)+1),
		E    => MODE,
		Q    => ConfigBits((k*2)+1) ); 
end generate;

CONFout <= ConfigBits(ConfigBits'high);  

--begin
--	if clk'event and CLK='1' then
--		if mode='1' then	--configuration mode
--		LUT_values <= LUT_values(LUT_values'high-1 downto 0) & CONFin;
--		c_out_mux  <= LUT_values(LUT_values'high);
--		c_I0mux    <= c_out_mux;
--		end if;
--	end if;
--end process;

LUT_values <= ConfigBits(15 downto 0);
c_out_mux  <= ConfigBits(16);
c_I0mux    <= ConfigBits(17);

--CONFout <= c_I0mux;

I0mux <= I0 when (c_I0mux = '0') else Ci;
LUT_index <= I3 & I2 & I1 & I0mux;

-- The LUT is just a multiplexer 
-- for a first shot, I am using a 16:1
-- LUT_out <= LUT_values(TO_INTEGER(LUT_index));
inst_MUX16PTv2_E6BEG1 : MUX16PTv2
	 Port Map(
		IN1 	=> LUT_values(0),
		IN2 	=> LUT_values(1),
		IN3 	=> LUT_values(2),
		IN4 	=> LUT_values(3),
		IN5 	=> LUT_values(4),
		IN6 	=> LUT_values(5),
		IN7 	=> LUT_values(6),
		IN8 	=> LUT_values(7),
		IN9 	=> LUT_values(8),
		IN10 	=> LUT_values(9),
		IN11 	=> LUT_values(10),
		IN12 	=> LUT_values(11),
		IN13 	=> LUT_values(12),
		IN14 	=> LUT_values(13),
		IN15 	=> LUT_values(14),
		IN16 	=> LUT_values(15),
		S1 	=> LUT_index(0),
		S2 	=> LUT_index(1),
		S3 	=> LUT_index(2),
		S4 	=> LUT_index(3),
		O  	=> LUT_out );

O <= LUT_flop when (c_out_mux = '1') else LUT_out;

Co <= (Ci AND I1) OR (Ci AND I2) OR (I1 AND I2);	-- iCE40 like carry chain (as this is supported in Josys; would normally go for fractured LUT

process(UserCLK)
begin
	if UserCLK'event and UserCLK='1' then
		LUT_flop <= LUT_out;
	end if;
end process;


end architecture Behavioral;
